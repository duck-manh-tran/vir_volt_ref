
.option MEASFORM=3
.param vdd=0.8
.param vinit=0.4

.ic v(vdis)='vinit+0.01'

.meas tran t_dis TRIG v(vdis) val='vinit' FALL=1 TARG v(vdis) val='vdd*0.25' FALL=1

.tran 1n 4m sweep DATA=input

.DATA input
+ vdd vinit
0.600 0.270
0.600 0.300
0.600 0.330
0.600 0.360
0.600 0.390
0.600 0.420
0.600 0.450
0.600 0.480
0.600 0.510
0.600 0.540
0.600 0.570
0.600 0.600
0.620 0.279
0.620 0.310
0.620 0.341
0.620 0.372
0.620 0.403
0.620 0.434
0.620 0.465
0.620 0.496
0.620 0.527
0.620 0.558
0.620 0.589
0.620 0.620
0.640 0.288
0.640 0.320
0.640 0.352
0.640 0.384
0.640 0.416
0.640 0.448
0.640 0.480
0.640 0.512
0.640 0.544
0.640 0.576
0.640 0.608
0.640 0.640
0.660 0.297
0.660 0.330
0.660 0.363
0.660 0.396
0.660 0.429
0.660 0.462
0.660 0.495
0.660 0.528
0.660 0.561
0.660 0.594
0.660 0.627
0.660 0.660
0.680 0.306
0.680 0.340
0.680 0.374
0.680 0.408
0.680 0.442
0.680 0.476
0.680 0.510
0.680 0.544
0.680 0.578
0.680 0.612
0.680 0.646
0.680 0.680
0.700 0.315
0.700 0.350
0.700 0.385
0.700 0.420
0.700 0.455
0.700 0.490
0.700 0.525
0.700 0.560
0.700 0.595
0.700 0.630
0.700 0.665
0.700 0.700
0.720 0.324
0.720 0.360
0.720 0.396
0.720 0.432
0.720 0.468
0.720 0.504
0.720 0.540
0.720 0.576
0.720 0.612
0.720 0.648
0.720 0.684
0.720 0.720
0.740 0.333
0.740 0.370
0.740 0.407
0.740 0.444
0.740 0.481
0.740 0.518
0.740 0.555
0.740 0.592
0.740 0.629
0.740 0.666
0.740 0.703
0.740 0.740
0.760 0.342
0.760 0.380
0.760 0.418
0.760 0.456
0.760 0.494
0.760 0.532
0.760 0.570
0.760 0.608
0.760 0.646
0.760 0.684
0.760 0.722
0.760 0.760
0.780 0.351
0.780 0.390
0.780 0.429
0.780 0.468
0.780 0.507
0.780 0.546
0.780 0.585
0.780 0.624
0.780 0.663
0.780 0.702
0.780 0.741
0.780 0.780
0.800 0.360
0.800 0.400
0.800 0.440
0.800 0.480
0.800 0.520
0.800 0.560
0.800 0.600
0.800 0.640
0.800 0.680
0.800 0.720
0.800 0.760
0.800 0.800
0.820 0.369
0.820 0.410
0.820 0.451
0.820 0.492
0.820 0.533
0.820 0.574
0.820 0.615
0.820 0.656
0.820 0.697
0.820 0.738
0.820 0.779
0.820 0.820
0.840 0.378
0.840 0.420
0.840 0.462
0.840 0.504
0.840 0.546
0.840 0.588
0.840 0.630
0.840 0.672
0.840 0.714
0.840 0.756
0.840 0.798
0.840 0.840
0.860 0.387
0.860 0.430
0.860 0.473
0.860 0.516
0.860 0.559
0.860 0.602
0.860 0.645
0.860 0.688
0.860 0.731
0.860 0.774
0.860 0.817
0.860 0.860
0.880 0.396
0.880 0.440
0.880 0.484
0.880 0.528
0.880 0.572
0.880 0.616
0.880 0.660
0.880 0.704
0.880 0.748
0.880 0.792
0.880 0.836
0.880 0.880
0.900 0.405
0.900 0.450
0.900 0.495
0.900 0.540
0.900 0.585
0.900 0.630
0.900 0.675
0.900 0.720
0.900 0.765
0.900 0.810
0.900 0.855
0.900 0.900
0.920 0.414
0.920 0.460
0.920 0.506
0.920 0.552
0.920 0.598
0.920 0.644
0.920 0.690
0.920 0.736
0.920 0.782
0.920 0.828
0.920 0.874
0.920 0.920
0.940 0.423
0.940 0.470
0.940 0.517
0.940 0.564
0.940 0.611
0.940 0.658
0.940 0.705
0.940 0.752
0.940 0.799
0.940 0.846
0.940 0.893
0.940 0.940
0.960 0.432
0.960 0.480
0.960 0.528
0.960 0.576
0.960 0.624
0.960 0.672
0.960 0.720
0.960 0.768
0.960 0.816
0.960 0.864
0.960 0.912
0.960 0.960
0.980 0.441
0.980 0.490
0.980 0.539
0.980 0.588
0.980 0.637
0.980 0.686
0.980 0.735
0.980 0.784
0.980 0.833
0.980 0.882
0.980 0.931
0.980 0.980
1.000 0.450
1.000 0.500
1.000 0.550
1.000 0.600
1.000 0.650
1.000 0.700
1.000 0.750
1.000 0.800
1.000 0.850
1.000 0.900
1.000 0.950
1.000 1.000
1.020 0.459
1.020 0.510
1.020 0.561
1.020 0.612
1.020 0.663
1.020 0.714
1.020 0.765
1.020 0.816
1.020 0.867
1.020 0.918
1.020 0.969
1.020 1.020
1.040 0.468
1.040 0.520
1.040 0.572
1.040 0.624
1.040 0.676
1.040 0.728
1.040 0.780
1.040 0.832
1.040 0.884
1.040 0.936
1.040 0.988
1.040 1.040
1.060 0.477
1.060 0.530
1.060 0.583
1.060 0.636
1.060 0.689
1.060 0.742
1.060 0.795
1.060 0.848
1.060 0.901
1.060 0.954
1.060 1.007
1.060 1.060
1.080 0.486
1.080 0.540
1.080 0.594
1.080 0.648
1.080 0.702
1.080 0.756
1.080 0.810
1.080 0.864
1.080 0.918
1.080 0.972
1.080 1.026
1.080 1.080
1.100 0.495
1.100 0.550
1.100 0.605
1.100 0.660
1.100 0.715
1.100 0.770
1.100 0.825
1.100 0.880
1.100 0.935
1.100 0.990
1.100 1.045
1.100 1.100
1.120 0.504
1.120 0.560
1.120 0.616
1.120 0.672
1.120 0.728
1.120 0.784
1.120 0.840
1.120 0.896
1.120 0.952
1.120 1.008
1.120 1.064
1.120 1.120
1.140 0.513
1.140 0.570
1.140 0.627
1.140 0.684
1.140 0.741
1.140 0.798
1.140 0.855
1.140 0.912
1.140 0.969
1.140 1.026
1.140 1.083
1.140 1.140
1.160 0.522
1.160 0.580
1.160 0.638
1.160 0.696
1.160 0.754
1.160 0.812
1.160 0.870
1.160 0.928
1.160 0.986
1.160 1.044
1.160 1.102
1.160 1.160
1.180 0.531
1.180 0.590
1.180 0.649
1.180 0.708
1.180 0.767
1.180 0.826
1.180 0.885
1.180 0.944
1.180 1.003
1.180 1.062
1.180 1.121
1.180 1.180
1.200 0.540
1.200 0.600
1.200 0.660
1.200 0.720
1.200 0.780
1.200 0.840
1.200 0.900
1.200 0.960
1.200 1.020
1.200 1.080
1.200 1.140
1.200 1.200
.ENDDATA
