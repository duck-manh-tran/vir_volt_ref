
.option MEASFORM=3
.param vdd=0.8
.param vinit=0.4
.param k1 = 0.4
.param k2 = 0.3
.param k3 = 0.25
.param v_cap1='vdd*r_cap*k1'
.param v_cap1='vdd*r_cap*k2'
.param v_cap1='vdd*r_cap*k3'

.ic v(vdis)='vdd+0.01'

.meas tran t_dis1 TRIG v(vdis) val='v_cap1' FALL=1 TARG v(vdis) val='vdd*0.25' FALL=1
.meas tran t_dis2 TRIG v(vdis) val='v_cap2' FALL=1 TARG v(vdis) val='vdd*0.25' FALL=1
.meas tran t_dis3 TRIG v(vdis) val='v_cap3' FALL=1 TARG v(vdis) val='vdd*0.25' FALL=1

.tran 1n 4m sweep DATA=input

.DATA input
+ vdd r_cap
.ENDDATA
