
.ic  v(vc)=0.3
.param collect_mode = 0
.option runlvl=6
.option opfile=1 split_dp=1
.option probe=1
.probe tran v(*) level=1
.probe tran v(vc) v(ctrl_dsn) v(ctrl_dsn_bar) v(vir_gnd)

.tran 1n 30m sweep DATA=input

.DATA input
+ vdd
+ 0.40
+ 0.41
+ 0.42
+ 0.43
+ 0.44
+ 0.45
+ 0.46
+ 0.47
+ 0.48
+ 0.49
+ 0.50
+ 0.51
+ 0.52
+ 0.53
+ 0.54
+ 0.55
+ 0.56
+ 0.57
+ 0.58
+ 0.59
+ 0.60
+ 0.61
+ 0.62
+ 0.63
+ 0.64
+ 0.65
+ 0.66
+ 0.67
+ 0.68
+ 0.69
+ 0.70
+ 0.71
+ 0.72
+ 0.73
+ 0.74
+ 0.75
+ 0.76
+ 0.77
+ 0.78
+ 0.79
+ 0.80
.ENDDATA
