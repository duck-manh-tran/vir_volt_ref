

.option MEASFORM=3
.param vdd=0.8
.param init=1.0
.param vinit='vdd*init'
.temp = temp_val

.ic v(vp)='vinit+0.01'

.meas tran t_dis TRIG v(vp) val='vinit' FALL=1 TARG v(vp) val='vdd*0.25' FALL=1

.tran 100p 3m sweep DATA=input

.DATA input
+ temp_val init
+ -40.0 0.3
+ -30.0 0.3
+ -20.0 0.3
+ -10.0 0.3
+ 0.0 0.3
+ 10.0 0.3
+ 20.0 0.3
+ 30.0 0.3
+ 40.0 0.3
+ 50.0 0.3
+ 60.0 0.3
+ 70.0 0.3
+ 80.0 0.3
+ 90.0 0.3
+ 100.0 0.3
+ -40.0 0.4
+ -30.0 0.4
+ -20.0 0.4
+ -10.0 0.4
+ 0.0 0.4
+ 10.0 0.4
+ 20.0 0.4
+ 30.0 0.4
+ 40.0 0.4
+ 50.0 0.4
+ 60.0 0.4
+ 70.0 0.4
+ 80.0 0.4
+ 90.0 0.4
+ 100.0 0.4
+ -40.0 0.5
+ -30.0 0.5
+ -20.0 0.5
+ -10.0 0.5
+ 0.0 0.5
+ 10.0 0.5
+ 20.0 0.5
+ 30.0 0.5
+ 40.0 0.5
+ 50.0 0.5
+ 60.0 0.5
+ 70.0 0.5
+ 80.0 0.5
+ 90.0 0.5
+ 100.0 0.5
+ -40.0 0.6
+ -30.0 0.6
+ -20.0 0.6
+ -10.0 0.6
+ 0.0 0.6
+ 10.0 0.6
+ 20.0 0.6
+ 30.0 0.6
+ 40.0 0.6
+ 50.0 0.6
+ 60.0 0.6
+ 70.0 0.6
+ 80.0 0.6
+ 90.0 0.6
+ 100.0 0.6
+ -40.0 0.7
+ -30.0 0.7
+ -20.0 0.7
+ -10.0 0.7
+ 0.0 0.7
+ 10.0 0.7
+ 20.0 0.7
+ 30.0 0.7
+ 40.0 0.7
+ 50.0 0.7
+ 60.0 0.7
+ 70.0 0.7
+ 80.0 0.7
+ 90.0 0.7
+ 100.0 0.7
+ -40.0 0.8
+ -30.0 0.8
+ -20.0 0.8
+ -10.0 0.8
+ 0.0 0.8
+ 10.0 0.8
+ 20.0 0.8
+ 30.0 0.8
+ 40.0 0.8
+ 50.0 0.8
+ 60.0 0.8
+ 70.0 0.8
+ 80.0 0.8
+ 90.0 0.8
+ 100.0 0.8
+ -40.0 0.9
+ -30.0 0.9
+ -20.0 0.9
+ -10.0 0.9
+ 0.0 0.9
+ 10.0 0.9
+ 20.0 0.9
+ 30.0 0.9
+ 40.0 0.9
+ 50.0 0.9
+ 60.0 0.9
+ 70.0 0.9
+ 80.0 0.9
+ 90.0 0.9
+ 100.0 0.9
+ -40.0 1.0
+ -30.0 1.0
+ -20.0 1.0
+ -10.0 1.0
+ 0.0 1.0
+ 10.0 1.0
+ 20.0 1.0
+ 30.0 1.0
+ 40.0 1.0
+ 50.0 1.0
+ 60.0 1.0
+ 70.0 1.0
+ 80.0 1.0
+ 90.0 1.0
+ 100.0 1.0
.ENDDATA
