
.option MEASFORM=3
.option RUNLVL=5
.option MEASDGT=6
.param vdd=0.8
.param vinit=0.4
.param k1 = 0.4
.param k2 = 0.3
.param k3 = 0.25
.param v_cap1='vdd*r_cap*k1'
.param v_cap2='vdd*r_cap*k2'
.param v_cap3='vdd*r_cap*k3'

.ic v(vdis)='vdd+0.01'

.meas tran t_dis1 TRIG v(vdis) val='v_cap1' FALL=1 TARG v(vdis) val='vdd*0.25' FALL=1
.meas tran t_dis2 TRIG v(vdis) val='v_cap2' FALL=1 TARG v(vdis) val='vdd*0.25' FALL=1
.meas tran t_dis3 TRIG v(vdis) val='v_cap3' FALL=1 TARG v(vdis) val='vdd*0.25' FALL=1

.tran 1n 4m sweep DATA=input

.DATA input
+ vdd r_cap
+ 0.400 1.250
+ 0.400 1.275
+ 0.400 1.300
+ 0.400 1.325
+ 0.400 1.350
+ 0.400 1.375
+ 0.400 1.400
+ 0.400 1.425
+ 0.400 1.450
+ 0.400 1.475
+ 0.400 1.500
+ 0.400 1.525
+ 0.400 1.550
+ 0.400 1.575
+ 0.400 1.600
+ 0.400 1.625
+ 0.400 1.650
+ 0.400 1.675
+ 0.400 1.700
+ 0.400 1.725
+ 0.400 1.750
+ 0.400 1.775
+ 0.400 1.800
+ 0.400 1.825
+ 0.400 1.850
+ 0.400 1.875
+ 0.400 1.900
+ 0.400 1.925
+ 0.400 1.950
+ 0.400 1.975
+ 0.400 2.000
+ 0.400 2.025
+ 0.400 2.050
+ 0.400 2.075
+ 0.400 2.100
+ 0.400 2.125
+ 0.400 2.150
+ 0.400 2.175
+ 0.400 2.200
+ 0.400 2.225
+ 0.400 2.250
+ 0.400 2.275
+ 0.400 2.300
+ 0.400 2.325
+ 0.400 2.350
+ 0.400 2.375
+ 0.400 2.400
+ 0.400 2.425
+ 0.400 2.450
+ 0.400 2.475
+ 0.400 2.500
+ 0.420 1.250
+ 0.420 1.275
+ 0.420 1.300
+ 0.420 1.325
+ 0.420 1.350
+ 0.420 1.375
+ 0.420 1.400
+ 0.420 1.425
+ 0.420 1.450
+ 0.420 1.475
+ 0.420 1.500
+ 0.420 1.525
+ 0.420 1.550
+ 0.420 1.575
+ 0.420 1.600
+ 0.420 1.625
+ 0.420 1.650
+ 0.420 1.675
+ 0.420 1.700
+ 0.420 1.725
+ 0.420 1.750
+ 0.420 1.775
+ 0.420 1.800
+ 0.420 1.825
+ 0.420 1.850
+ 0.420 1.875
+ 0.420 1.900
+ 0.420 1.925
+ 0.420 1.950
+ 0.420 1.975
+ 0.420 2.000
+ 0.420 2.025
+ 0.420 2.050
+ 0.420 2.075
+ 0.420 2.100
+ 0.420 2.125
+ 0.420 2.150
+ 0.420 2.175
+ 0.420 2.200
+ 0.420 2.225
+ 0.420 2.250
+ 0.420 2.275
+ 0.420 2.300
+ 0.420 2.325
+ 0.420 2.350
+ 0.420 2.375
+ 0.420 2.400
+ 0.420 2.425
+ 0.420 2.450
+ 0.420 2.475
+ 0.420 2.500
+ 0.440 1.250
+ 0.440 1.275
+ 0.440 1.300
+ 0.440 1.325
+ 0.440 1.350
+ 0.440 1.375
+ 0.440 1.400
+ 0.440 1.425
+ 0.440 1.450
+ 0.440 1.475
+ 0.440 1.500
+ 0.440 1.525
+ 0.440 1.550
+ 0.440 1.575
+ 0.440 1.600
+ 0.440 1.625
+ 0.440 1.650
+ 0.440 1.675
+ 0.440 1.700
+ 0.440 1.725
+ 0.440 1.750
+ 0.440 1.775
+ 0.440 1.800
+ 0.440 1.825
+ 0.440 1.850
+ 0.440 1.875
+ 0.440 1.900
+ 0.440 1.925
+ 0.440 1.950
+ 0.440 1.975
+ 0.440 2.000
+ 0.440 2.025
+ 0.440 2.050
+ 0.440 2.075
+ 0.440 2.100
+ 0.440 2.125
+ 0.440 2.150
+ 0.440 2.175
+ 0.440 2.200
+ 0.440 2.225
+ 0.440 2.250
+ 0.440 2.275
+ 0.440 2.300
+ 0.440 2.325
+ 0.440 2.350
+ 0.440 2.375
+ 0.440 2.400
+ 0.440 2.425
+ 0.440 2.450
+ 0.440 2.475
+ 0.440 2.500
+ 0.460 1.250
+ 0.460 1.275
+ 0.460 1.300
+ 0.460 1.325
+ 0.460 1.350
+ 0.460 1.375
+ 0.460 1.400
+ 0.460 1.425
+ 0.460 1.450
+ 0.460 1.475
+ 0.460 1.500
+ 0.460 1.525
+ 0.460 1.550
+ 0.460 1.575
+ 0.460 1.600
+ 0.460 1.625
+ 0.460 1.650
+ 0.460 1.675
+ 0.460 1.700
+ 0.460 1.725
+ 0.460 1.750
+ 0.460 1.775
+ 0.460 1.800
+ 0.460 1.825
+ 0.460 1.850
+ 0.460 1.875
+ 0.460 1.900
+ 0.460 1.925
+ 0.460 1.950
+ 0.460 1.975
+ 0.460 2.000
+ 0.460 2.025
+ 0.460 2.050
+ 0.460 2.075
+ 0.460 2.100
+ 0.460 2.125
+ 0.460 2.150
+ 0.460 2.175
+ 0.460 2.200
+ 0.460 2.225
+ 0.460 2.250
+ 0.460 2.275
+ 0.460 2.300
+ 0.460 2.325
+ 0.460 2.350
+ 0.460 2.375
+ 0.460 2.400
+ 0.460 2.425
+ 0.460 2.450
+ 0.460 2.475
+ 0.460 2.500
+ 0.480 1.250
+ 0.480 1.275
+ 0.480 1.300
+ 0.480 1.325
+ 0.480 1.350
+ 0.480 1.375
+ 0.480 1.400
+ 0.480 1.425
+ 0.480 1.450
+ 0.480 1.475
+ 0.480 1.500
+ 0.480 1.525
+ 0.480 1.550
+ 0.480 1.575
+ 0.480 1.600
+ 0.480 1.625
+ 0.480 1.650
+ 0.480 1.675
+ 0.480 1.700
+ 0.480 1.725
+ 0.480 1.750
+ 0.480 1.775
+ 0.480 1.800
+ 0.480 1.825
+ 0.480 1.850
+ 0.480 1.875
+ 0.480 1.900
+ 0.480 1.925
+ 0.480 1.950
+ 0.480 1.975
+ 0.480 2.000
+ 0.480 2.025
+ 0.480 2.050
+ 0.480 2.075
+ 0.480 2.100
+ 0.480 2.125
+ 0.480 2.150
+ 0.480 2.175
+ 0.480 2.200
+ 0.480 2.225
+ 0.480 2.250
+ 0.480 2.275
+ 0.480 2.300
+ 0.480 2.325
+ 0.480 2.350
+ 0.480 2.375
+ 0.480 2.400
+ 0.480 2.425
+ 0.480 2.450
+ 0.480 2.475
+ 0.480 2.500
+ 0.500 1.250
+ 0.500 1.275
+ 0.500 1.300
+ 0.500 1.325
+ 0.500 1.350
+ 0.500 1.375
+ 0.500 1.400
+ 0.500 1.425
+ 0.500 1.450
+ 0.500 1.475
+ 0.500 1.500
+ 0.500 1.525
+ 0.500 1.550
+ 0.500 1.575
+ 0.500 1.600
+ 0.500 1.625
+ 0.500 1.650
+ 0.500 1.675
+ 0.500 1.700
+ 0.500 1.725
+ 0.500 1.750
+ 0.500 1.775
+ 0.500 1.800
+ 0.500 1.825
+ 0.500 1.850
+ 0.500 1.875
+ 0.500 1.900
+ 0.500 1.925
+ 0.500 1.950
+ 0.500 1.975
+ 0.500 2.000
+ 0.500 2.025
+ 0.500 2.050
+ 0.500 2.075
+ 0.500 2.100
+ 0.500 2.125
+ 0.500 2.150
+ 0.500 2.175
+ 0.500 2.200
+ 0.500 2.225
+ 0.500 2.250
+ 0.500 2.275
+ 0.500 2.300
+ 0.500 2.325
+ 0.500 2.350
+ 0.500 2.375
+ 0.500 2.400
+ 0.500 2.425
+ 0.500 2.450
+ 0.500 2.475
+ 0.500 2.500
+ 0.520 1.250
+ 0.520 1.275
+ 0.520 1.300
+ 0.520 1.325
+ 0.520 1.350
+ 0.520 1.375
+ 0.520 1.400
+ 0.520 1.425
+ 0.520 1.450
+ 0.520 1.475
+ 0.520 1.500
+ 0.520 1.525
+ 0.520 1.550
+ 0.520 1.575
+ 0.520 1.600
+ 0.520 1.625
+ 0.520 1.650
+ 0.520 1.675
+ 0.520 1.700
+ 0.520 1.725
+ 0.520 1.750
+ 0.520 1.775
+ 0.520 1.800
+ 0.520 1.825
+ 0.520 1.850
+ 0.520 1.875
+ 0.520 1.900
+ 0.520 1.925
+ 0.520 1.950
+ 0.520 1.975
+ 0.520 2.000
+ 0.520 2.025
+ 0.520 2.050
+ 0.520 2.075
+ 0.520 2.100
+ 0.520 2.125
+ 0.520 2.150
+ 0.520 2.175
+ 0.520 2.200
+ 0.520 2.225
+ 0.520 2.250
+ 0.520 2.275
+ 0.520 2.300
+ 0.520 2.325
+ 0.520 2.350
+ 0.520 2.375
+ 0.520 2.400
+ 0.520 2.425
+ 0.520 2.450
+ 0.520 2.475
+ 0.520 2.500
+ 0.540 1.250
+ 0.540 1.275
+ 0.540 1.300
+ 0.540 1.325
+ 0.540 1.350
+ 0.540 1.375
+ 0.540 1.400
+ 0.540 1.425
+ 0.540 1.450
+ 0.540 1.475
+ 0.540 1.500
+ 0.540 1.525
+ 0.540 1.550
+ 0.540 1.575
+ 0.540 1.600
+ 0.540 1.625
+ 0.540 1.650
+ 0.540 1.675
+ 0.540 1.700
+ 0.540 1.725
+ 0.540 1.750
+ 0.540 1.775
+ 0.540 1.800
+ 0.540 1.825
+ 0.540 1.850
+ 0.540 1.875
+ 0.540 1.900
+ 0.540 1.925
+ 0.540 1.950
+ 0.540 1.975
+ 0.540 2.000
+ 0.540 2.025
+ 0.540 2.050
+ 0.540 2.075
+ 0.540 2.100
+ 0.540 2.125
+ 0.540 2.150
+ 0.540 2.175
+ 0.540 2.200
+ 0.540 2.225
+ 0.540 2.250
+ 0.540 2.275
+ 0.540 2.300
+ 0.540 2.325
+ 0.540 2.350
+ 0.540 2.375
+ 0.540 2.400
+ 0.540 2.425
+ 0.540 2.450
+ 0.540 2.475
+ 0.540 2.500
+ 0.560 1.250
+ 0.560 1.275
+ 0.560 1.300
+ 0.560 1.325
+ 0.560 1.350
+ 0.560 1.375
+ 0.560 1.400
+ 0.560 1.425
+ 0.560 1.450
+ 0.560 1.475
+ 0.560 1.500
+ 0.560 1.525
+ 0.560 1.550
+ 0.560 1.575
+ 0.560 1.600
+ 0.560 1.625
+ 0.560 1.650
+ 0.560 1.675
+ 0.560 1.700
+ 0.560 1.725
+ 0.560 1.750
+ 0.560 1.775
+ 0.560 1.800
+ 0.560 1.825
+ 0.560 1.850
+ 0.560 1.875
+ 0.560 1.900
+ 0.560 1.925
+ 0.560 1.950
+ 0.560 1.975
+ 0.560 2.000
+ 0.560 2.025
+ 0.560 2.050
+ 0.560 2.075
+ 0.560 2.100
+ 0.560 2.125
+ 0.560 2.150
+ 0.560 2.175
+ 0.560 2.200
+ 0.560 2.225
+ 0.560 2.250
+ 0.560 2.275
+ 0.560 2.300
+ 0.560 2.325
+ 0.560 2.350
+ 0.560 2.375
+ 0.560 2.400
+ 0.560 2.425
+ 0.560 2.450
+ 0.560 2.475
+ 0.560 2.500
+ 0.580 1.250
+ 0.580 1.275
+ 0.580 1.300
+ 0.580 1.325
+ 0.580 1.350
+ 0.580 1.375
+ 0.580 1.400
+ 0.580 1.425
+ 0.580 1.450
+ 0.580 1.475
+ 0.580 1.500
+ 0.580 1.525
+ 0.580 1.550
+ 0.580 1.575
+ 0.580 1.600
+ 0.580 1.625
+ 0.580 1.650
+ 0.580 1.675
+ 0.580 1.700
+ 0.580 1.725
+ 0.580 1.750
+ 0.580 1.775
+ 0.580 1.800
+ 0.580 1.825
+ 0.580 1.850
+ 0.580 1.875
+ 0.580 1.900
+ 0.580 1.925
+ 0.580 1.950
+ 0.580 1.975
+ 0.580 2.000
+ 0.580 2.025
+ 0.580 2.050
+ 0.580 2.075
+ 0.580 2.100
+ 0.580 2.125
+ 0.580 2.150
+ 0.580 2.175
+ 0.580 2.200
+ 0.580 2.225
+ 0.580 2.250
+ 0.580 2.275
+ 0.580 2.300
+ 0.580 2.325
+ 0.580 2.350
+ 0.580 2.375
+ 0.580 2.400
+ 0.580 2.425
+ 0.580 2.450
+ 0.580 2.475
+ 0.580 2.500
+ 0.600 1.250
+ 0.600 1.275
+ 0.600 1.300
+ 0.600 1.325
+ 0.600 1.350
+ 0.600 1.375
+ 0.600 1.400
+ 0.600 1.425
+ 0.600 1.450
+ 0.600 1.475
+ 0.600 1.500
+ 0.600 1.525
+ 0.600 1.550
+ 0.600 1.575
+ 0.600 1.600
+ 0.600 1.625
+ 0.600 1.650
+ 0.600 1.675
+ 0.600 1.700
+ 0.600 1.725
+ 0.600 1.750
+ 0.600 1.775
+ 0.600 1.800
+ 0.600 1.825
+ 0.600 1.850
+ 0.600 1.875
+ 0.600 1.900
+ 0.600 1.925
+ 0.600 1.950
+ 0.600 1.975
+ 0.600 2.000
+ 0.600 2.025
+ 0.600 2.050
+ 0.600 2.075
+ 0.600 2.100
+ 0.600 2.125
+ 0.600 2.150
+ 0.600 2.175
+ 0.600 2.200
+ 0.600 2.225
+ 0.600 2.250
+ 0.600 2.275
+ 0.600 2.300
+ 0.600 2.325
+ 0.600 2.350
+ 0.600 2.375
+ 0.600 2.400
+ 0.600 2.425
+ 0.600 2.450
+ 0.600 2.475
+ 0.600 2.500
+ 0.620 1.250
+ 0.620 1.275
+ 0.620 1.300
+ 0.620 1.325
+ 0.620 1.350
+ 0.620 1.375
+ 0.620 1.400
+ 0.620 1.425
+ 0.620 1.450
+ 0.620 1.475
+ 0.620 1.500
+ 0.620 1.525
+ 0.620 1.550
+ 0.620 1.575
+ 0.620 1.600
+ 0.620 1.625
+ 0.620 1.650
+ 0.620 1.675
+ 0.620 1.700
+ 0.620 1.725
+ 0.620 1.750
+ 0.620 1.775
+ 0.620 1.800
+ 0.620 1.825
+ 0.620 1.850
+ 0.620 1.875
+ 0.620 1.900
+ 0.620 1.925
+ 0.620 1.950
+ 0.620 1.975
+ 0.620 2.000
+ 0.620 2.025
+ 0.620 2.050
+ 0.620 2.075
+ 0.620 2.100
+ 0.620 2.125
+ 0.620 2.150
+ 0.620 2.175
+ 0.620 2.200
+ 0.620 2.225
+ 0.620 2.250
+ 0.620 2.275
+ 0.620 2.300
+ 0.620 2.325
+ 0.620 2.350
+ 0.620 2.375
+ 0.620 2.400
+ 0.620 2.425
+ 0.620 2.450
+ 0.620 2.475
+ 0.620 2.500
+ 0.640 1.250
+ 0.640 1.275
+ 0.640 1.300
+ 0.640 1.325
+ 0.640 1.350
+ 0.640 1.375
+ 0.640 1.400
+ 0.640 1.425
+ 0.640 1.450
+ 0.640 1.475
+ 0.640 1.500
+ 0.640 1.525
+ 0.640 1.550
+ 0.640 1.575
+ 0.640 1.600
+ 0.640 1.625
+ 0.640 1.650
+ 0.640 1.675
+ 0.640 1.700
+ 0.640 1.725
+ 0.640 1.750
+ 0.640 1.775
+ 0.640 1.800
+ 0.640 1.825
+ 0.640 1.850
+ 0.640 1.875
+ 0.640 1.900
+ 0.640 1.925
+ 0.640 1.950
+ 0.640 1.975
+ 0.640 2.000
+ 0.640 2.025
+ 0.640 2.050
+ 0.640 2.075
+ 0.640 2.100
+ 0.640 2.125
+ 0.640 2.150
+ 0.640 2.175
+ 0.640 2.200
+ 0.640 2.225
+ 0.640 2.250
+ 0.640 2.275
+ 0.640 2.300
+ 0.640 2.325
+ 0.640 2.350
+ 0.640 2.375
+ 0.640 2.400
+ 0.640 2.425
+ 0.640 2.450
+ 0.640 2.475
+ 0.640 2.500
+ 0.660 1.250
+ 0.660 1.275
+ 0.660 1.300
+ 0.660 1.325
+ 0.660 1.350
+ 0.660 1.375
+ 0.660 1.400
+ 0.660 1.425
+ 0.660 1.450
+ 0.660 1.475
+ 0.660 1.500
+ 0.660 1.525
+ 0.660 1.550
+ 0.660 1.575
+ 0.660 1.600
+ 0.660 1.625
+ 0.660 1.650
+ 0.660 1.675
+ 0.660 1.700
+ 0.660 1.725
+ 0.660 1.750
+ 0.660 1.775
+ 0.660 1.800
+ 0.660 1.825
+ 0.660 1.850
+ 0.660 1.875
+ 0.660 1.900
+ 0.660 1.925
+ 0.660 1.950
+ 0.660 1.975
+ 0.660 2.000
+ 0.660 2.025
+ 0.660 2.050
+ 0.660 2.075
+ 0.660 2.100
+ 0.660 2.125
+ 0.660 2.150
+ 0.660 2.175
+ 0.660 2.200
+ 0.660 2.225
+ 0.660 2.250
+ 0.660 2.275
+ 0.660 2.300
+ 0.660 2.325
+ 0.660 2.350
+ 0.660 2.375
+ 0.660 2.400
+ 0.660 2.425
+ 0.660 2.450
+ 0.660 2.475
+ 0.660 2.500
+ 0.680 1.250
+ 0.680 1.275
+ 0.680 1.300
+ 0.680 1.325
+ 0.680 1.350
+ 0.680 1.375
+ 0.680 1.400
+ 0.680 1.425
+ 0.680 1.450
+ 0.680 1.475
+ 0.680 1.500
+ 0.680 1.525
+ 0.680 1.550
+ 0.680 1.575
+ 0.680 1.600
+ 0.680 1.625
+ 0.680 1.650
+ 0.680 1.675
+ 0.680 1.700
+ 0.680 1.725
+ 0.680 1.750
+ 0.680 1.775
+ 0.680 1.800
+ 0.680 1.825
+ 0.680 1.850
+ 0.680 1.875
+ 0.680 1.900
+ 0.680 1.925
+ 0.680 1.950
+ 0.680 1.975
+ 0.680 2.000
+ 0.680 2.025
+ 0.680 2.050
+ 0.680 2.075
+ 0.680 2.100
+ 0.680 2.125
+ 0.680 2.150
+ 0.680 2.175
+ 0.680 2.200
+ 0.680 2.225
+ 0.680 2.250
+ 0.680 2.275
+ 0.680 2.300
+ 0.680 2.325
+ 0.680 2.350
+ 0.680 2.375
+ 0.680 2.400
+ 0.680 2.425
+ 0.680 2.450
+ 0.680 2.475
+ 0.680 2.500
+ 0.700 1.250
+ 0.700 1.275
+ 0.700 1.300
+ 0.700 1.325
+ 0.700 1.350
+ 0.700 1.375
+ 0.700 1.400
+ 0.700 1.425
+ 0.700 1.450
+ 0.700 1.475
+ 0.700 1.500
+ 0.700 1.525
+ 0.700 1.550
+ 0.700 1.575
+ 0.700 1.600
+ 0.700 1.625
+ 0.700 1.650
+ 0.700 1.675
+ 0.700 1.700
+ 0.700 1.725
+ 0.700 1.750
+ 0.700 1.775
+ 0.700 1.800
+ 0.700 1.825
+ 0.700 1.850
+ 0.700 1.875
+ 0.700 1.900
+ 0.700 1.925
+ 0.700 1.950
+ 0.700 1.975
+ 0.700 2.000
+ 0.700 2.025
+ 0.700 2.050
+ 0.700 2.075
+ 0.700 2.100
+ 0.700 2.125
+ 0.700 2.150
+ 0.700 2.175
+ 0.700 2.200
+ 0.700 2.225
+ 0.700 2.250
+ 0.700 2.275
+ 0.700 2.300
+ 0.700 2.325
+ 0.700 2.350
+ 0.700 2.375
+ 0.700 2.400
+ 0.700 2.425
+ 0.700 2.450
+ 0.700 2.475
+ 0.700 2.500
+ 0.720 1.250
+ 0.720 1.275
+ 0.720 1.300
+ 0.720 1.325
+ 0.720 1.350
+ 0.720 1.375
+ 0.720 1.400
+ 0.720 1.425
+ 0.720 1.450
+ 0.720 1.475
+ 0.720 1.500
+ 0.720 1.525
+ 0.720 1.550
+ 0.720 1.575
+ 0.720 1.600
+ 0.720 1.625
+ 0.720 1.650
+ 0.720 1.675
+ 0.720 1.700
+ 0.720 1.725
+ 0.720 1.750
+ 0.720 1.775
+ 0.720 1.800
+ 0.720 1.825
+ 0.720 1.850
+ 0.720 1.875
+ 0.720 1.900
+ 0.720 1.925
+ 0.720 1.950
+ 0.720 1.975
+ 0.720 2.000
+ 0.720 2.025
+ 0.720 2.050
+ 0.720 2.075
+ 0.720 2.100
+ 0.720 2.125
+ 0.720 2.150
+ 0.720 2.175
+ 0.720 2.200
+ 0.720 2.225
+ 0.720 2.250
+ 0.720 2.275
+ 0.720 2.300
+ 0.720 2.325
+ 0.720 2.350
+ 0.720 2.375
+ 0.720 2.400
+ 0.720 2.425
+ 0.720 2.450
+ 0.720 2.475
+ 0.720 2.500
+ 0.740 1.250
+ 0.740 1.275
+ 0.740 1.300
+ 0.740 1.325
+ 0.740 1.350
+ 0.740 1.375
+ 0.740 1.400
+ 0.740 1.425
+ 0.740 1.450
+ 0.740 1.475
+ 0.740 1.500
+ 0.740 1.525
+ 0.740 1.550
+ 0.740 1.575
+ 0.740 1.600
+ 0.740 1.625
+ 0.740 1.650
+ 0.740 1.675
+ 0.740 1.700
+ 0.740 1.725
+ 0.740 1.750
+ 0.740 1.775
+ 0.740 1.800
+ 0.740 1.825
+ 0.740 1.850
+ 0.740 1.875
+ 0.740 1.900
+ 0.740 1.925
+ 0.740 1.950
+ 0.740 1.975
+ 0.740 2.000
+ 0.740 2.025
+ 0.740 2.050
+ 0.740 2.075
+ 0.740 2.100
+ 0.740 2.125
+ 0.740 2.150
+ 0.740 2.175
+ 0.740 2.200
+ 0.740 2.225
+ 0.740 2.250
+ 0.740 2.275
+ 0.740 2.300
+ 0.740 2.325
+ 0.740 2.350
+ 0.740 2.375
+ 0.740 2.400
+ 0.740 2.425
+ 0.740 2.450
+ 0.740 2.475
+ 0.740 2.500
+ 0.760 1.250
+ 0.760 1.275
+ 0.760 1.300
+ 0.760 1.325
+ 0.760 1.350
+ 0.760 1.375
+ 0.760 1.400
+ 0.760 1.425
+ 0.760 1.450
+ 0.760 1.475
+ 0.760 1.500
+ 0.760 1.525
+ 0.760 1.550
+ 0.760 1.575
+ 0.760 1.600
+ 0.760 1.625
+ 0.760 1.650
+ 0.760 1.675
+ 0.760 1.700
+ 0.760 1.725
+ 0.760 1.750
+ 0.760 1.775
+ 0.760 1.800
+ 0.760 1.825
+ 0.760 1.850
+ 0.760 1.875
+ 0.760 1.900
+ 0.760 1.925
+ 0.760 1.950
+ 0.760 1.975
+ 0.760 2.000
+ 0.760 2.025
+ 0.760 2.050
+ 0.760 2.075
+ 0.760 2.100
+ 0.760 2.125
+ 0.760 2.150
+ 0.760 2.175
+ 0.760 2.200
+ 0.760 2.225
+ 0.760 2.250
+ 0.760 2.275
+ 0.760 2.300
+ 0.760 2.325
+ 0.760 2.350
+ 0.760 2.375
+ 0.760 2.400
+ 0.760 2.425
+ 0.760 2.450
+ 0.760 2.475
+ 0.760 2.500
+ 0.780 1.250
+ 0.780 1.275
+ 0.780 1.300
+ 0.780 1.325
+ 0.780 1.350
+ 0.780 1.375
+ 0.780 1.400
+ 0.780 1.425
+ 0.780 1.450
+ 0.780 1.475
+ 0.780 1.500
+ 0.780 1.525
+ 0.780 1.550
+ 0.780 1.575
+ 0.780 1.600
+ 0.780 1.625
+ 0.780 1.650
+ 0.780 1.675
+ 0.780 1.700
+ 0.780 1.725
+ 0.780 1.750
+ 0.780 1.775
+ 0.780 1.800
+ 0.780 1.825
+ 0.780 1.850
+ 0.780 1.875
+ 0.780 1.900
+ 0.780 1.925
+ 0.780 1.950
+ 0.780 1.975
+ 0.780 2.000
+ 0.780 2.025
+ 0.780 2.050
+ 0.780 2.075
+ 0.780 2.100
+ 0.780 2.125
+ 0.780 2.150
+ 0.780 2.175
+ 0.780 2.200
+ 0.780 2.225
+ 0.780 2.250
+ 0.780 2.275
+ 0.780 2.300
+ 0.780 2.325
+ 0.780 2.350
+ 0.780 2.375
+ 0.780 2.400
+ 0.780 2.425
+ 0.780 2.450
+ 0.780 2.475
+ 0.780 2.500
+ 0.800 1.250
+ 0.800 1.275
+ 0.800 1.300
+ 0.800 1.325
+ 0.800 1.350
+ 0.800 1.375
+ 0.800 1.400
+ 0.800 1.425
+ 0.800 1.450
+ 0.800 1.475
+ 0.800 1.500
+ 0.800 1.525
+ 0.800 1.550
+ 0.800 1.575
+ 0.800 1.600
+ 0.800 1.625
+ 0.800 1.650
+ 0.800 1.675
+ 0.800 1.700
+ 0.800 1.725
+ 0.800 1.750
+ 0.800 1.775
+ 0.800 1.800
+ 0.800 1.825
+ 0.800 1.850
+ 0.800 1.875
+ 0.800 1.900
+ 0.800 1.925
+ 0.800 1.950
+ 0.800 1.975
+ 0.800 2.000
+ 0.800 2.025
+ 0.800 2.050
+ 0.800 2.075
+ 0.800 2.100
+ 0.800 2.125
+ 0.800 2.150
+ 0.800 2.175
+ 0.800 2.200
+ 0.800 2.225
+ 0.800 2.250
+ 0.800 2.275
+ 0.800 2.300
+ 0.800 2.325
+ 0.800 2.350
+ 0.800 2.375
+ 0.800 2.400
+ 0.800 2.425
+ 0.800 2.450
+ 0.800 2.475
+ 0.800 2.500
.ENDDATA
