** circuit: digital_BGR_model

.subckt discharge_nwk _VP_ VGND W=0.5
XM1 net3 net3 _VP_ _VP_ sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM2 net2 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM3 net1 net1 net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1 
XM4 net4 net4 net2 net2 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM5 GND VGND net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XC1 _VP_ VGND sky130_fd_pr__cap_mim_m3_2 W=14.5 L=1.5 MF=10 m=10
.ends

X_discharge_nwk VP GND discharge_nwk W=W
 
* Digital circuits by xspice
a8 enb %gd(VP_ VP) switch3
.model switch3 aswitch(cntl_off=0.0 cntl_on=0.4 r_off=1e15
+ r_on=10k log=TRUE limit=TRUE)

* Voltage setup for the circuit
V_DAC VP_ GND DC=0.05
V_sup VDD GND DC=v_dd
V_enb enb GND pulse (0 v_dd T_set 0 0 T_on 1 1)
V_clk clk GND pulse (0 0.8 0 'prd/20' 'prd/20' '9*prd/20' prd)

* Setup simulation 
.lib ~/work/conda_eda/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.param clk_freq = 1e6
.param prd = '1/clk_freq'
.param T_set = 0.1m T_on = 0.5m
.param W = 0.5
.param V_init = 0.2
.param v_dd = 0.8
.csparam v_dd_ = {v_dd}
.ic v(VP) = V_init
.option trtol = 5

.control
save all
echo  ______________________________________
echo |   go to the measurement operation    |
echo  --------------------------------------
let NoL = 65536		$ Number of DAC Levels
let m = vector(3)		$ storage of DAC m levels
let n = vector(3)		$ storage of TDC discharge time
let DAC_vol = vector(3)		$ storage of the DAC voltage
* get the value of the m vector
let ix = 0
while (ix<3)
	let m[ix] = `/bin/bash -c "python processor_model.py $&ix"`
	let DAC_vol[ix] = (m[ix]/NoL)*v_dd_
	let ix = ix+1
end

stop when v(enb) > 0.4  when v(VP_) = 0.05

let quad_dvol1 = DAC_vol[0]/4
let dvol1 = DAC_vol[0]-0.01
stop when v(VP)<'$&quad_dvol1' when v(VP_) ge '$&dvol1'

let quad_dvol2 = DAC_vol[1]/4
let dvol2 = DAC_vol[1]-0.01
stop when v(VP)<'$&quad_dvol2' when v(VP_) ge '$&dvol2'

* let quad_dvol3 = DAC_vol[2]/4
* let dvol3 = DAC_vol[2]-0.01
* stop when v(VP)<'$&quad_dvol3' when v(VP_) ge '$&dvol3'

tran 100n 80m

alter V_DAC dc = DAC_vol[0]
resume

meas tran t1_stop when v(VP) = '$&quad_dvol1' CROSS=1
let t1_charge = t1_stop+0.1m
alter @V_enb[pulse] = (0 '$&v_dd_' '$&t1_charge' 0 0 0.5m 1)
alter V_DAC dc = DAC_vol[1]
resume

meas tran t2_stop when v(VP) = '$&quad_dvol2' CROSS=1
let t2_charge = t2_stop+0.1m
alter @V_enb[pulse] = (0 '$&v_dd_' '$&t2_charge' 0 0 0.5m 1)
alter V_DAC dc = DAC_vol[2]
resume


plot enb vp vp_
.endc
**** end user architecture code
**.ends
.GLOBAL GND
.end

* alter V_DAC dc=DAC_vol
* alter V_sup dc=$v_dd
* let quad_dd = $v_dd/4
* meas tran DAC_out AVG v(VP_) from=2m to=10m
* meas tran t_dis WHEN v(VP)=quad_dd CROSS=LAST
* meas tran t_dis trig v(enb) val=0 FALL=1  targ v(VP) val=quad_dd FALL=1
* let n[im] = 't_dis-1.1m'
* print DAC_out
* let im = im+1
* end
* print n > discharge_time.txt
* write d_bgr_model.raw
* 
* echo " _________________________________________"
* echo "|   go to the reference hold operation		|"
* echo " -----------------------------------------"
* 
* save VP_ VP enb clk  
* set N = 65536
* let DAC_vol = ($m_set/$N)*$v_dd
* alter V_sup dc=$v_dd
* alter V_DAC dc=DAC_vol
* run
* let ix=ix+1
* meas tran DAC_out AVG v(VP_) from=2m to=10m
* print DAC_out
* end
* write d_bgr_model.raw
* 

