** sch_path: /home/manhtd_61d/work/d_bgr/xschem/discharge_nwk.sch
**.subckt discharge_nwk

.subckt discharge_nwk ctrl VP VGND W=0.5 L=0.15
** diode based transistors
XM1 net1 net1 VP 	VP	 sky130_fd_pr__pfet_01v8 L="L" W=W nf=1 
XM2 net2 net2 net1 net1 sky130_fd_pr__pfet_01v8 L="L" W=W nf=1 
XM3 net3 net3 net2 net2 sky130_fd_pr__pfet_01v8 L="L" W=W nf=1 
XM4 net4 net4 net3 net3 sky130_fd_pr__pfet_01v8 L="L" W=W nf=1 
XM5 net5 net5 net4 net4 sky130_fd_pr__pfet_01v8 L="L" W=W nf=1 
XML netk netk net5 net5 sky130_fd_pr__pfet_01v8 L="L" W=W nf=1 
** locker
Xk1 netk ctrl VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=2 
Xk2 netk ctrl VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=2 
Xsky130_fd_pr__cap_vpp0 VP VGND VGND VGND sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 m=1
Xsky130_fd_pr__cap_vpp1 VP VGND VGND VGND sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 m=1
Xsky130_fd_pr__cap_vpp2 VP VGND VGND VGND sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 m=1
Xsky130_fd_pr__cap_vpp3 VP VGND VGND VGND sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 m=1
.ends

.subckt discharge_nwk1 ctrl _VP_ VGND W=0.5
XM1 net3 net3 _VP_ _VP_ sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM2 net2 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM3 net1 net1 net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM4 net4 net4 net2 net2 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM5 netk netk net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
Xsky130_fd_pr__cap_vpp0 _VP_ VGND VGND VGND sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 m=1
Xsky130_fd_pr__cap_vpp1 _VP_ VGND VGND VGND sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 m=1
Xsky130_fd_pr__cap_vpp2 _VP_ VGND VGND VGND sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 m=1
Xsky130_fd_pr__cap_vpp3 _VP_ VGND VGND VGND sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 m=1
XMk netk ctrl VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=2
.ends

X_discharge_nwk ctrl VP1 GND discharge_nwk W=W L=L
* X_discharge_nwk1 ctrl VP1 GND discharge_nwk1 W=W
**** begin user architecture code

.lib /home/dkits/efabless/mpw-7a/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice hh
.param W = 1
.param L = 0.18
.param V_init = 0.81
.param v_dd = 0.8
*.ic v(VP0) = V_init
.ic v(VP1) = V_init

V_ctrl ctrl gnd dc='v_dd'
* V_DAC res_net gnd dc='v_dd'
* R1 res_net VP1 r = 10000
.control
set num_threads=12
save VP1 ctrl

set temp = $temp_c
tran $step_time $stop_time

print VP1 > ./result/temp/l180nm/nf_6/$outfile
quit

.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
