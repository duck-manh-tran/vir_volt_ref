
.ic  v(vc)=0.3
.param collect_mode = 0
.option runlvl=6
.option opfile=1 split_dp=1
.option probe=1
.probe tran v(*) level=1
.probe tran v(vc) v(ctrl_dsn) v(ctrl_dsn_bar) v(vir_gnd)

.tran 1n 30m sweep DATA=input

.DATA input
+ vdd r_cap
+ 0.4 1.25
+ 0.4 1.26
+ 0.4 1.27
+ 0.4 1.28
+ 0.4 1.29
+ 0.4 1.3
+ 0.4 1.31
+ 0.4 1.32
+ 0.4 1.33
+ 0.4 1.34
+ 0.4 1.35
+ 0.4 1.36
+ 0.4 1.37
+ 0.4 1.38
+ 0.4 1.39
+ 0.4 1.4
+ 0.4 1.41
+ 0.4 1.42
+ 0.4 1.43
+ 0.4 1.44
+ 0.4 1.45
+ 0.4 1.46
+ 0.4 1.47
+ 0.4 1.48
+ 0.4 1.49
+ 0.4 1.5
+ 0.4 1.51
+ 0.4 1.52
+ 0.4 1.53
+ 0.4 1.54
+ 0.4 1.55
+ 0.4 1.56
+ 0.4 1.57
+ 0.4 1.58
+ 0.4 1.59
+ 0.4 1.6
+ 0.4 1.61
+ 0.4 1.62
+ 0.4 1.63
+ 0.4 1.64
+ 0.4 1.65
+ 0.4 1.66
+ 0.4 1.67
+ 0.4 1.68
+ 0.4 1.69
+ 0.4 1.7
+ 0.4 1.71
+ 0.4 1.72
+ 0.4 1.73
+ 0.4 1.74
+ 0.4 1.75
+ 0.4 1.76
+ 0.4 1.77
+ 0.4 1.78
+ 0.4 1.79
+ 0.4 1.8
+ 0.4 1.81
+ 0.4 1.82
+ 0.4 1.83
+ 0.4 1.84
+ 0.4 1.85
+ 0.4 1.86
+ 0.4 1.87
+ 0.4 1.88
+ 0.4 1.89
+ 0.4 1.9
+ 0.4 1.91
+ 0.4 1.92
+ 0.4 1.93
+ 0.4 1.94
+ 0.4 1.95
+ 0.4 1.96
+ 0.4 1.97
+ 0.4 1.98
+ 0.4 1.99
+ 0.4 2.0
+ 0.4 2.01
+ 0.4 2.02
+ 0.4 2.03
+ 0.4 2.04
+ 0.4 2.05
+ 0.4 2.06
+ 0.4 2.07
+ 0.4 2.08
+ 0.4 2.09
+ 0.4 2.1
+ 0.4 2.11
+ 0.4 2.12
+ 0.4 2.13
+ 0.4 2.14
+ 0.4 2.15
+ 0.4 2.16
+ 0.4 2.17
+ 0.4 2.18
+ 0.4 2.19
+ 0.4 2.2
+ 0.4 2.21
+ 0.4 2.22
+ 0.4 2.23
+ 0.4 2.24
+ 0.4 2.25
+ 0.4 2.26
+ 0.4 2.27
+ 0.4 2.28
+ 0.4 2.29
+ 0.4 2.3
+ 0.4 2.31
+ 0.4 2.32
+ 0.4 2.33
+ 0.4 2.34
+ 0.4 2.35
+ 0.4 2.36
+ 0.4 2.37
+ 0.4 2.38
+ 0.4 2.39
+ 0.4 2.4
+ 0.4 2.41
+ 0.4 2.42
+ 0.4 2.43
+ 0.4 2.44
+ 0.4 2.45
+ 0.4 2.46
+ 0.4 2.47
+ 0.4 2.48
+ 0.4 2.49
+ 0.4 2.5
+ 0.41 1.25
+ 0.41 1.26
+ 0.41 1.27
+ 0.41 1.28
+ 0.41 1.29
+ 0.41 1.3
+ 0.41 1.31
+ 0.41 1.32
+ 0.41 1.33
+ 0.41 1.34
+ 0.41 1.35
+ 0.41 1.36
+ 0.41 1.37
+ 0.41 1.38
+ 0.41 1.39
+ 0.41 1.4
+ 0.41 1.41
+ 0.41 1.42
+ 0.41 1.43
+ 0.41 1.44
+ 0.41 1.45
+ 0.41 1.46
+ 0.41 1.47
+ 0.41 1.48
+ 0.41 1.49
+ 0.41 1.5
+ 0.41 1.51
+ 0.41 1.52
+ 0.41 1.53
+ 0.41 1.54
+ 0.41 1.55
+ 0.41 1.56
+ 0.41 1.57
+ 0.41 1.58
+ 0.41 1.59
+ 0.41 1.6
+ 0.41 1.61
+ 0.41 1.62
+ 0.41 1.63
+ 0.41 1.64
+ 0.41 1.65
+ 0.41 1.66
+ 0.41 1.67
+ 0.41 1.68
+ 0.41 1.69
+ 0.41 1.7
+ 0.41 1.71
+ 0.41 1.72
+ 0.41 1.73
+ 0.41 1.74
+ 0.41 1.75
+ 0.41 1.76
+ 0.41 1.77
+ 0.41 1.78
+ 0.41 1.79
+ 0.41 1.8
+ 0.41 1.81
+ 0.41 1.82
+ 0.41 1.83
+ 0.41 1.84
+ 0.41 1.85
+ 0.41 1.86
+ 0.41 1.87
+ 0.41 1.88
+ 0.41 1.89
+ 0.41 1.9
+ 0.41 1.91
+ 0.41 1.92
+ 0.41 1.93
+ 0.41 1.94
+ 0.41 1.95
+ 0.41 1.96
+ 0.41 1.97
+ 0.41 1.98
+ 0.41 1.99
+ 0.41 2.0
+ 0.41 2.01
+ 0.41 2.02
+ 0.41 2.03
+ 0.41 2.04
+ 0.41 2.05
+ 0.41 2.06
+ 0.41 2.07
+ 0.41 2.08
+ 0.41 2.09
+ 0.41 2.1
+ 0.41 2.11
+ 0.41 2.12
+ 0.41 2.13
+ 0.41 2.14
+ 0.41 2.15
+ 0.41 2.16
+ 0.41 2.17
+ 0.41 2.18
+ 0.41 2.19
+ 0.41 2.2
+ 0.41 2.21
+ 0.41 2.22
+ 0.41 2.23
+ 0.41 2.24
+ 0.41 2.25
+ 0.41 2.26
+ 0.41 2.27
+ 0.41 2.28
+ 0.41 2.29
+ 0.41 2.3
+ 0.41 2.31
+ 0.41 2.32
+ 0.41 2.33
+ 0.41 2.34
+ 0.41 2.35
+ 0.41 2.36
+ 0.41 2.37
+ 0.41 2.38
+ 0.41 2.39
+ 0.41 2.4
+ 0.41 2.41
+ 0.41 2.42
+ 0.41 2.43
+ 0.41 2.44
+ 0.41 2.45
+ 0.41 2.46
+ 0.41 2.47
+ 0.41 2.48
+ 0.41 2.49
+ 0.41 2.5
+ 0.42 1.25
+ 0.42 1.26
+ 0.42 1.27
+ 0.42 1.28
+ 0.42 1.29
+ 0.42 1.3
+ 0.42 1.31
+ 0.42 1.32
+ 0.42 1.33
+ 0.42 1.34
+ 0.42 1.35
+ 0.42 1.36
+ 0.42 1.37
+ 0.42 1.38
+ 0.42 1.39
+ 0.42 1.4
+ 0.42 1.41
+ 0.42 1.42
+ 0.42 1.43
+ 0.42 1.44
+ 0.42 1.45
+ 0.42 1.46
+ 0.42 1.47
+ 0.42 1.48
+ 0.42 1.49
+ 0.42 1.5
+ 0.42 1.51
+ 0.42 1.52
+ 0.42 1.53
+ 0.42 1.54
+ 0.42 1.55
+ 0.42 1.56
+ 0.42 1.57
+ 0.42 1.58
+ 0.42 1.59
+ 0.42 1.6
+ 0.42 1.61
+ 0.42 1.62
+ 0.42 1.63
+ 0.42 1.64
+ 0.42 1.65
+ 0.42 1.66
+ 0.42 1.67
+ 0.42 1.68
+ 0.42 1.69
+ 0.42 1.7
+ 0.42 1.71
+ 0.42 1.72
+ 0.42 1.73
+ 0.42 1.74
+ 0.42 1.75
+ 0.42 1.76
+ 0.42 1.77
+ 0.42 1.78
+ 0.42 1.79
+ 0.42 1.8
+ 0.42 1.81
+ 0.42 1.82
+ 0.42 1.83
+ 0.42 1.84
+ 0.42 1.85
+ 0.42 1.86
+ 0.42 1.87
+ 0.42 1.88
+ 0.42 1.89
+ 0.42 1.9
+ 0.42 1.91
+ 0.42 1.92
+ 0.42 1.93
+ 0.42 1.94
+ 0.42 1.95
+ 0.42 1.96
+ 0.42 1.97
+ 0.42 1.98
+ 0.42 1.99
+ 0.42 2.0
+ 0.42 2.01
+ 0.42 2.02
+ 0.42 2.03
+ 0.42 2.04
+ 0.42 2.05
+ 0.42 2.06
+ 0.42 2.07
+ 0.42 2.08
+ 0.42 2.09
+ 0.42 2.1
+ 0.42 2.11
+ 0.42 2.12
+ 0.42 2.13
+ 0.42 2.14
+ 0.42 2.15
+ 0.42 2.16
+ 0.42 2.17
+ 0.42 2.18
+ 0.42 2.19
+ 0.42 2.2
+ 0.42 2.21
+ 0.42 2.22
+ 0.42 2.23
+ 0.42 2.24
+ 0.42 2.25
+ 0.42 2.26
+ 0.42 2.27
+ 0.42 2.28
+ 0.42 2.29
+ 0.42 2.3
+ 0.42 2.31
+ 0.42 2.32
+ 0.42 2.33
+ 0.42 2.34
+ 0.42 2.35
+ 0.42 2.36
+ 0.42 2.37
+ 0.42 2.38
+ 0.42 2.39
+ 0.42 2.4
+ 0.42 2.41
+ 0.42 2.42
+ 0.42 2.43
+ 0.42 2.44
+ 0.42 2.45
+ 0.42 2.46
+ 0.42 2.47
+ 0.42 2.48
+ 0.42 2.49
+ 0.42 2.5
+ 0.43 1.25
+ 0.43 1.26
+ 0.43 1.27
+ 0.43 1.28
+ 0.43 1.29
+ 0.43 1.3
+ 0.43 1.31
+ 0.43 1.32
+ 0.43 1.33
+ 0.43 1.34
+ 0.43 1.35
+ 0.43 1.36
+ 0.43 1.37
+ 0.43 1.38
+ 0.43 1.39
+ 0.43 1.4
+ 0.43 1.41
+ 0.43 1.42
+ 0.43 1.43
+ 0.43 1.44
+ 0.43 1.45
+ 0.43 1.46
+ 0.43 1.47
+ 0.43 1.48
+ 0.43 1.49
+ 0.43 1.5
+ 0.43 1.51
+ 0.43 1.52
+ 0.43 1.53
+ 0.43 1.54
+ 0.43 1.55
+ 0.43 1.56
+ 0.43 1.57
+ 0.43 1.58
+ 0.43 1.59
+ 0.43 1.6
+ 0.43 1.61
+ 0.43 1.62
+ 0.43 1.63
+ 0.43 1.64
+ 0.43 1.65
+ 0.43 1.66
+ 0.43 1.67
+ 0.43 1.68
+ 0.43 1.69
+ 0.43 1.7
+ 0.43 1.71
+ 0.43 1.72
+ 0.43 1.73
+ 0.43 1.74
+ 0.43 1.75
+ 0.43 1.76
+ 0.43 1.77
+ 0.43 1.78
+ 0.43 1.79
+ 0.43 1.8
+ 0.43 1.81
+ 0.43 1.82
+ 0.43 1.83
+ 0.43 1.84
+ 0.43 1.85
+ 0.43 1.86
+ 0.43 1.87
+ 0.43 1.88
+ 0.43 1.89
+ 0.43 1.9
+ 0.43 1.91
+ 0.43 1.92
+ 0.43 1.93
+ 0.43 1.94
+ 0.43 1.95
+ 0.43 1.96
+ 0.43 1.97
+ 0.43 1.98
+ 0.43 1.99
+ 0.43 2.0
+ 0.43 2.01
+ 0.43 2.02
+ 0.43 2.03
+ 0.43 2.04
+ 0.43 2.05
+ 0.43 2.06
+ 0.43 2.07
+ 0.43 2.08
+ 0.43 2.09
+ 0.43 2.1
+ 0.43 2.11
+ 0.43 2.12
+ 0.43 2.13
+ 0.43 2.14
+ 0.43 2.15
+ 0.43 2.16
+ 0.43 2.17
+ 0.43 2.18
+ 0.43 2.19
+ 0.43 2.2
+ 0.43 2.21
+ 0.43 2.22
+ 0.43 2.23
+ 0.43 2.24
+ 0.43 2.25
+ 0.43 2.26
+ 0.43 2.27
+ 0.43 2.28
+ 0.43 2.29
+ 0.43 2.3
+ 0.43 2.31
+ 0.43 2.32
+ 0.43 2.33
+ 0.43 2.34
+ 0.43 2.35
+ 0.43 2.36
+ 0.43 2.37
+ 0.43 2.38
+ 0.43 2.39
+ 0.43 2.4
+ 0.43 2.41
+ 0.43 2.42
+ 0.43 2.43
+ 0.43 2.44
+ 0.43 2.45
+ 0.43 2.46
+ 0.43 2.47
+ 0.43 2.48
+ 0.43 2.49
+ 0.43 2.5
+ 0.44 1.25
+ 0.44 1.26
+ 0.44 1.27
+ 0.44 1.28
+ 0.44 1.29
+ 0.44 1.3
+ 0.44 1.31
+ 0.44 1.32
+ 0.44 1.33
+ 0.44 1.34
+ 0.44 1.35
+ 0.44 1.36
+ 0.44 1.37
+ 0.44 1.38
+ 0.44 1.39
+ 0.44 1.4
+ 0.44 1.41
+ 0.44 1.42
+ 0.44 1.43
+ 0.44 1.44
+ 0.44 1.45
+ 0.44 1.46
+ 0.44 1.47
+ 0.44 1.48
+ 0.44 1.49
+ 0.44 1.5
+ 0.44 1.51
+ 0.44 1.52
+ 0.44 1.53
+ 0.44 1.54
+ 0.44 1.55
+ 0.44 1.56
+ 0.44 1.57
+ 0.44 1.58
+ 0.44 1.59
+ 0.44 1.6
+ 0.44 1.61
+ 0.44 1.62
+ 0.44 1.63
+ 0.44 1.64
+ 0.44 1.65
+ 0.44 1.66
+ 0.44 1.67
+ 0.44 1.68
+ 0.44 1.69
+ 0.44 1.7
+ 0.44 1.71
+ 0.44 1.72
+ 0.44 1.73
+ 0.44 1.74
+ 0.44 1.75
+ 0.44 1.76
+ 0.44 1.77
+ 0.44 1.78
+ 0.44 1.79
+ 0.44 1.8
+ 0.44 1.81
+ 0.44 1.82
+ 0.44 1.83
+ 0.44 1.84
+ 0.44 1.85
+ 0.44 1.86
+ 0.44 1.87
+ 0.44 1.88
+ 0.44 1.89
+ 0.44 1.9
+ 0.44 1.91
+ 0.44 1.92
+ 0.44 1.93
+ 0.44 1.94
+ 0.44 1.95
+ 0.44 1.96
+ 0.44 1.97
+ 0.44 1.98
+ 0.44 1.99
+ 0.44 2.0
+ 0.44 2.01
+ 0.44 2.02
+ 0.44 2.03
+ 0.44 2.04
+ 0.44 2.05
+ 0.44 2.06
+ 0.44 2.07
+ 0.44 2.08
+ 0.44 2.09
+ 0.44 2.1
+ 0.44 2.11
+ 0.44 2.12
+ 0.44 2.13
+ 0.44 2.14
+ 0.44 2.15
+ 0.44 2.16
+ 0.44 2.17
+ 0.44 2.18
+ 0.44 2.19
+ 0.44 2.2
+ 0.44 2.21
+ 0.44 2.22
+ 0.44 2.23
+ 0.44 2.24
+ 0.44 2.25
+ 0.44 2.26
+ 0.44 2.27
+ 0.44 2.28
+ 0.44 2.29
+ 0.44 2.3
+ 0.44 2.31
+ 0.44 2.32
+ 0.44 2.33
+ 0.44 2.34
+ 0.44 2.35
+ 0.44 2.36
+ 0.44 2.37
+ 0.44 2.38
+ 0.44 2.39
+ 0.44 2.4
+ 0.44 2.41
+ 0.44 2.42
+ 0.44 2.43
+ 0.44 2.44
+ 0.44 2.45
+ 0.44 2.46
+ 0.44 2.47
+ 0.44 2.48
+ 0.44 2.49
+ 0.44 2.5
+ 0.45 1.25
+ 0.45 1.26
+ 0.45 1.27
+ 0.45 1.28
+ 0.45 1.29
+ 0.45 1.3
+ 0.45 1.31
+ 0.45 1.32
+ 0.45 1.33
+ 0.45 1.34
+ 0.45 1.35
+ 0.45 1.36
+ 0.45 1.37
+ 0.45 1.38
+ 0.45 1.39
+ 0.45 1.4
+ 0.45 1.41
+ 0.45 1.42
+ 0.45 1.43
+ 0.45 1.44
+ 0.45 1.45
+ 0.45 1.46
+ 0.45 1.47
+ 0.45 1.48
+ 0.45 1.49
+ 0.45 1.5
+ 0.45 1.51
+ 0.45 1.52
+ 0.45 1.53
+ 0.45 1.54
+ 0.45 1.55
+ 0.45 1.56
+ 0.45 1.57
+ 0.45 1.58
+ 0.45 1.59
+ 0.45 1.6
+ 0.45 1.61
+ 0.45 1.62
+ 0.45 1.63
+ 0.45 1.64
+ 0.45 1.65
+ 0.45 1.66
+ 0.45 1.67
+ 0.45 1.68
+ 0.45 1.69
+ 0.45 1.7
+ 0.45 1.71
+ 0.45 1.72
+ 0.45 1.73
+ 0.45 1.74
+ 0.45 1.75
+ 0.45 1.76
+ 0.45 1.77
+ 0.45 1.78
+ 0.45 1.79
+ 0.45 1.8
+ 0.45 1.81
+ 0.45 1.82
+ 0.45 1.83
+ 0.45 1.84
+ 0.45 1.85
+ 0.45 1.86
+ 0.45 1.87
+ 0.45 1.88
+ 0.45 1.89
+ 0.45 1.9
+ 0.45 1.91
+ 0.45 1.92
+ 0.45 1.93
+ 0.45 1.94
+ 0.45 1.95
+ 0.45 1.96
+ 0.45 1.97
+ 0.45 1.98
+ 0.45 1.99
+ 0.45 2.0
+ 0.45 2.01
+ 0.45 2.02
+ 0.45 2.03
+ 0.45 2.04
+ 0.45 2.05
+ 0.45 2.06
+ 0.45 2.07
+ 0.45 2.08
+ 0.45 2.09
+ 0.45 2.1
+ 0.45 2.11
+ 0.45 2.12
+ 0.45 2.13
+ 0.45 2.14
+ 0.45 2.15
+ 0.45 2.16
+ 0.45 2.17
+ 0.45 2.18
+ 0.45 2.19
+ 0.45 2.2
+ 0.45 2.21
+ 0.45 2.22
+ 0.45 2.23
+ 0.45 2.24
+ 0.45 2.25
+ 0.45 2.26
+ 0.45 2.27
+ 0.45 2.28
+ 0.45 2.29
+ 0.45 2.3
+ 0.45 2.31
+ 0.45 2.32
+ 0.45 2.33
+ 0.45 2.34
+ 0.45 2.35
+ 0.45 2.36
+ 0.45 2.37
+ 0.45 2.38
+ 0.45 2.39
+ 0.45 2.4
+ 0.45 2.41
+ 0.45 2.42
+ 0.45 2.43
+ 0.45 2.44
+ 0.45 2.45
+ 0.45 2.46
+ 0.45 2.47
+ 0.45 2.48
+ 0.45 2.49
+ 0.45 2.5
+ 0.46 1.25
+ 0.46 1.26
+ 0.46 1.27
+ 0.46 1.28
+ 0.46 1.29
+ 0.46 1.3
+ 0.46 1.31
+ 0.46 1.32
+ 0.46 1.33
+ 0.46 1.34
+ 0.46 1.35
+ 0.46 1.36
+ 0.46 1.37
+ 0.46 1.38
+ 0.46 1.39
+ 0.46 1.4
+ 0.46 1.41
+ 0.46 1.42
+ 0.46 1.43
+ 0.46 1.44
+ 0.46 1.45
+ 0.46 1.46
+ 0.46 1.47
+ 0.46 1.48
+ 0.46 1.49
+ 0.46 1.5
+ 0.46 1.51
+ 0.46 1.52
+ 0.46 1.53
+ 0.46 1.54
+ 0.46 1.55
+ 0.46 1.56
+ 0.46 1.57
+ 0.46 1.58
+ 0.46 1.59
+ 0.46 1.6
+ 0.46 1.61
+ 0.46 1.62
+ 0.46 1.63
+ 0.46 1.64
+ 0.46 1.65
+ 0.46 1.66
+ 0.46 1.67
+ 0.46 1.68
+ 0.46 1.69
+ 0.46 1.7
+ 0.46 1.71
+ 0.46 1.72
+ 0.46 1.73
+ 0.46 1.74
+ 0.46 1.75
+ 0.46 1.76
+ 0.46 1.77
+ 0.46 1.78
+ 0.46 1.79
+ 0.46 1.8
+ 0.46 1.81
+ 0.46 1.82
+ 0.46 1.83
+ 0.46 1.84
+ 0.46 1.85
+ 0.46 1.86
+ 0.46 1.87
+ 0.46 1.88
+ 0.46 1.89
+ 0.46 1.9
+ 0.46 1.91
+ 0.46 1.92
+ 0.46 1.93
+ 0.46 1.94
+ 0.46 1.95
+ 0.46 1.96
+ 0.46 1.97
+ 0.46 1.98
+ 0.46 1.99
+ 0.46 2.0
+ 0.46 2.01
+ 0.46 2.02
+ 0.46 2.03
+ 0.46 2.04
+ 0.46 2.05
+ 0.46 2.06
+ 0.46 2.07
+ 0.46 2.08
+ 0.46 2.09
+ 0.46 2.1
+ 0.46 2.11
+ 0.46 2.12
+ 0.46 2.13
+ 0.46 2.14
+ 0.46 2.15
+ 0.46 2.16
+ 0.46 2.17
+ 0.46 2.18
+ 0.46 2.19
+ 0.46 2.2
+ 0.46 2.21
+ 0.46 2.22
+ 0.46 2.23
+ 0.46 2.24
+ 0.46 2.25
+ 0.46 2.26
+ 0.46 2.27
+ 0.46 2.28
+ 0.46 2.29
+ 0.46 2.3
+ 0.46 2.31
+ 0.46 2.32
+ 0.46 2.33
+ 0.46 2.34
+ 0.46 2.35
+ 0.46 2.36
+ 0.46 2.37
+ 0.46 2.38
+ 0.46 2.39
+ 0.46 2.4
+ 0.46 2.41
+ 0.46 2.42
+ 0.46 2.43
+ 0.46 2.44
+ 0.46 2.45
+ 0.46 2.46
+ 0.46 2.47
+ 0.46 2.48
+ 0.46 2.49
+ 0.46 2.5
+ 0.47 1.25
+ 0.47 1.26
+ 0.47 1.27
+ 0.47 1.28
+ 0.47 1.29
+ 0.47 1.3
+ 0.47 1.31
+ 0.47 1.32
+ 0.47 1.33
+ 0.47 1.34
+ 0.47 1.35
+ 0.47 1.36
+ 0.47 1.37
+ 0.47 1.38
+ 0.47 1.39
+ 0.47 1.4
+ 0.47 1.41
+ 0.47 1.42
+ 0.47 1.43
+ 0.47 1.44
+ 0.47 1.45
+ 0.47 1.46
+ 0.47 1.47
+ 0.47 1.48
+ 0.47 1.49
+ 0.47 1.5
+ 0.47 1.51
+ 0.47 1.52
+ 0.47 1.53
+ 0.47 1.54
+ 0.47 1.55
+ 0.47 1.56
+ 0.47 1.57
+ 0.47 1.58
+ 0.47 1.59
+ 0.47 1.6
+ 0.47 1.61
+ 0.47 1.62
+ 0.47 1.63
+ 0.47 1.64
+ 0.47 1.65
+ 0.47 1.66
+ 0.47 1.67
+ 0.47 1.68
+ 0.47 1.69
+ 0.47 1.7
+ 0.47 1.71
+ 0.47 1.72
+ 0.47 1.73
+ 0.47 1.74
+ 0.47 1.75
+ 0.47 1.76
+ 0.47 1.77
+ 0.47 1.78
+ 0.47 1.79
+ 0.47 1.8
+ 0.47 1.81
+ 0.47 1.82
+ 0.47 1.83
+ 0.47 1.84
+ 0.47 1.85
+ 0.47 1.86
+ 0.47 1.87
+ 0.47 1.88
+ 0.47 1.89
+ 0.47 1.9
+ 0.47 1.91
+ 0.47 1.92
+ 0.47 1.93
+ 0.47 1.94
+ 0.47 1.95
+ 0.47 1.96
+ 0.47 1.97
+ 0.47 1.98
+ 0.47 1.99
+ 0.47 2.0
+ 0.47 2.01
+ 0.47 2.02
+ 0.47 2.03
+ 0.47 2.04
+ 0.47 2.05
+ 0.47 2.06
+ 0.47 2.07
+ 0.47 2.08
+ 0.47 2.09
+ 0.47 2.1
+ 0.47 2.11
+ 0.47 2.12
+ 0.47 2.13
+ 0.47 2.14
+ 0.47 2.15
+ 0.47 2.16
+ 0.47 2.17
+ 0.47 2.18
+ 0.47 2.19
+ 0.47 2.2
+ 0.47 2.21
+ 0.47 2.22
+ 0.47 2.23
+ 0.47 2.24
+ 0.47 2.25
+ 0.47 2.26
+ 0.47 2.27
+ 0.47 2.28
+ 0.47 2.29
+ 0.47 2.3
+ 0.47 2.31
+ 0.47 2.32
+ 0.47 2.33
+ 0.47 2.34
+ 0.47 2.35
+ 0.47 2.36
+ 0.47 2.37
+ 0.47 2.38
+ 0.47 2.39
+ 0.47 2.4
+ 0.47 2.41
+ 0.47 2.42
+ 0.47 2.43
+ 0.47 2.44
+ 0.47 2.45
+ 0.47 2.46
+ 0.47 2.47
+ 0.47 2.48
+ 0.47 2.49
+ 0.47 2.5
+ 0.48 1.25
+ 0.48 1.26
+ 0.48 1.27
+ 0.48 1.28
+ 0.48 1.29
+ 0.48 1.3
+ 0.48 1.31
+ 0.48 1.32
+ 0.48 1.33
+ 0.48 1.34
+ 0.48 1.35
+ 0.48 1.36
+ 0.48 1.37
+ 0.48 1.38
+ 0.48 1.39
+ 0.48 1.4
+ 0.48 1.41
+ 0.48 1.42
+ 0.48 1.43
+ 0.48 1.44
+ 0.48 1.45
+ 0.48 1.46
+ 0.48 1.47
+ 0.48 1.48
+ 0.48 1.49
+ 0.48 1.5
+ 0.48 1.51
+ 0.48 1.52
+ 0.48 1.53
+ 0.48 1.54
+ 0.48 1.55
+ 0.48 1.56
+ 0.48 1.57
+ 0.48 1.58
+ 0.48 1.59
+ 0.48 1.6
+ 0.48 1.61
+ 0.48 1.62
+ 0.48 1.63
+ 0.48 1.64
+ 0.48 1.65
+ 0.48 1.66
+ 0.48 1.67
+ 0.48 1.68
+ 0.48 1.69
+ 0.48 1.7
+ 0.48 1.71
+ 0.48 1.72
+ 0.48 1.73
+ 0.48 1.74
+ 0.48 1.75
+ 0.48 1.76
+ 0.48 1.77
+ 0.48 1.78
+ 0.48 1.79
+ 0.48 1.8
+ 0.48 1.81
+ 0.48 1.82
+ 0.48 1.83
+ 0.48 1.84
+ 0.48 1.85
+ 0.48 1.86
+ 0.48 1.87
+ 0.48 1.88
+ 0.48 1.89
+ 0.48 1.9
+ 0.48 1.91
+ 0.48 1.92
+ 0.48 1.93
+ 0.48 1.94
+ 0.48 1.95
+ 0.48 1.96
+ 0.48 1.97
+ 0.48 1.98
+ 0.48 1.99
+ 0.48 2.0
+ 0.48 2.01
+ 0.48 2.02
+ 0.48 2.03
+ 0.48 2.04
+ 0.48 2.05
+ 0.48 2.06
+ 0.48 2.07
+ 0.48 2.08
+ 0.48 2.09
+ 0.48 2.1
+ 0.48 2.11
+ 0.48 2.12
+ 0.48 2.13
+ 0.48 2.14
+ 0.48 2.15
+ 0.48 2.16
+ 0.48 2.17
+ 0.48 2.18
+ 0.48 2.19
+ 0.48 2.2
+ 0.48 2.21
+ 0.48 2.22
+ 0.48 2.23
+ 0.48 2.24
+ 0.48 2.25
+ 0.48 2.26
+ 0.48 2.27
+ 0.48 2.28
+ 0.48 2.29
+ 0.48 2.3
+ 0.48 2.31
+ 0.48 2.32
+ 0.48 2.33
+ 0.48 2.34
+ 0.48 2.35
+ 0.48 2.36
+ 0.48 2.37
+ 0.48 2.38
+ 0.48 2.39
+ 0.48 2.4
+ 0.48 2.41
+ 0.48 2.42
+ 0.48 2.43
+ 0.48 2.44
+ 0.48 2.45
+ 0.48 2.46
+ 0.48 2.47
+ 0.48 2.48
+ 0.48 2.49
+ 0.48 2.5
+ 0.49 1.25
+ 0.49 1.26
+ 0.49 1.27
+ 0.49 1.28
+ 0.49 1.29
+ 0.49 1.3
+ 0.49 1.31
+ 0.49 1.32
+ 0.49 1.33
+ 0.49 1.34
+ 0.49 1.35
+ 0.49 1.36
+ 0.49 1.37
+ 0.49 1.38
+ 0.49 1.39
+ 0.49 1.4
+ 0.49 1.41
+ 0.49 1.42
+ 0.49 1.43
+ 0.49 1.44
+ 0.49 1.45
+ 0.49 1.46
+ 0.49 1.47
+ 0.49 1.48
+ 0.49 1.49
+ 0.49 1.5
+ 0.49 1.51
+ 0.49 1.52
+ 0.49 1.53
+ 0.49 1.54
+ 0.49 1.55
+ 0.49 1.56
+ 0.49 1.57
+ 0.49 1.58
+ 0.49 1.59
+ 0.49 1.6
+ 0.49 1.61
+ 0.49 1.62
+ 0.49 1.63
+ 0.49 1.64
+ 0.49 1.65
+ 0.49 1.66
+ 0.49 1.67
+ 0.49 1.68
+ 0.49 1.69
+ 0.49 1.7
+ 0.49 1.71
+ 0.49 1.72
+ 0.49 1.73
+ 0.49 1.74
+ 0.49 1.75
+ 0.49 1.76
+ 0.49 1.77
+ 0.49 1.78
+ 0.49 1.79
+ 0.49 1.8
+ 0.49 1.81
+ 0.49 1.82
+ 0.49 1.83
+ 0.49 1.84
+ 0.49 1.85
+ 0.49 1.86
+ 0.49 1.87
+ 0.49 1.88
+ 0.49 1.89
+ 0.49 1.9
+ 0.49 1.91
+ 0.49 1.92
+ 0.49 1.93
+ 0.49 1.94
+ 0.49 1.95
+ 0.49 1.96
+ 0.49 1.97
+ 0.49 1.98
+ 0.49 1.99
+ 0.49 2.0
+ 0.49 2.01
+ 0.49 2.02
+ 0.49 2.03
+ 0.49 2.04
+ 0.49 2.05
+ 0.49 2.06
+ 0.49 2.07
+ 0.49 2.08
+ 0.49 2.09
+ 0.49 2.1
+ 0.49 2.11
+ 0.49 2.12
+ 0.49 2.13
+ 0.49 2.14
+ 0.49 2.15
+ 0.49 2.16
+ 0.49 2.17
+ 0.49 2.18
+ 0.49 2.19
+ 0.49 2.2
+ 0.49 2.21
+ 0.49 2.22
+ 0.49 2.23
+ 0.49 2.24
+ 0.49 2.25
+ 0.49 2.26
+ 0.49 2.27
+ 0.49 2.28
+ 0.49 2.29
+ 0.49 2.3
+ 0.49 2.31
+ 0.49 2.32
+ 0.49 2.33
+ 0.49 2.34
+ 0.49 2.35
+ 0.49 2.36
+ 0.49 2.37
+ 0.49 2.38
+ 0.49 2.39
+ 0.49 2.4
+ 0.49 2.41
+ 0.49 2.42
+ 0.49 2.43
+ 0.49 2.44
+ 0.49 2.45
+ 0.49 2.46
+ 0.49 2.47
+ 0.49 2.48
+ 0.49 2.49
+ 0.49 2.5
+ 0.5 1.25
+ 0.5 1.26
+ 0.5 1.27
+ 0.5 1.28
+ 0.5 1.29
+ 0.5 1.3
+ 0.5 1.31
+ 0.5 1.32
+ 0.5 1.33
+ 0.5 1.34
+ 0.5 1.35
+ 0.5 1.36
+ 0.5 1.37
+ 0.5 1.38
+ 0.5 1.39
+ 0.5 1.4
+ 0.5 1.41
+ 0.5 1.42
+ 0.5 1.43
+ 0.5 1.44
+ 0.5 1.45
+ 0.5 1.46
+ 0.5 1.47
+ 0.5 1.48
+ 0.5 1.49
+ 0.5 1.5
+ 0.5 1.51
+ 0.5 1.52
+ 0.5 1.53
+ 0.5 1.54
+ 0.5 1.55
+ 0.5 1.56
+ 0.5 1.57
+ 0.5 1.58
+ 0.5 1.59
+ 0.5 1.6
+ 0.5 1.61
+ 0.5 1.62
+ 0.5 1.63
+ 0.5 1.64
+ 0.5 1.65
+ 0.5 1.66
+ 0.5 1.67
+ 0.5 1.68
+ 0.5 1.69
+ 0.5 1.7
+ 0.5 1.71
+ 0.5 1.72
+ 0.5 1.73
+ 0.5 1.74
+ 0.5 1.75
+ 0.5 1.76
+ 0.5 1.77
+ 0.5 1.78
+ 0.5 1.79
+ 0.5 1.8
+ 0.5 1.81
+ 0.5 1.82
+ 0.5 1.83
+ 0.5 1.84
+ 0.5 1.85
+ 0.5 1.86
+ 0.5 1.87
+ 0.5 1.88
+ 0.5 1.89
+ 0.5 1.9
+ 0.5 1.91
+ 0.5 1.92
+ 0.5 1.93
+ 0.5 1.94
+ 0.5 1.95
+ 0.5 1.96
+ 0.5 1.97
+ 0.5 1.98
+ 0.5 1.99
+ 0.5 2.0
+ 0.5 2.01
+ 0.5 2.02
+ 0.5 2.03
+ 0.5 2.04
+ 0.5 2.05
+ 0.5 2.06
+ 0.5 2.07
+ 0.5 2.08
+ 0.5 2.09
+ 0.5 2.1
+ 0.5 2.11
+ 0.5 2.12
+ 0.5 2.13
+ 0.5 2.14
+ 0.5 2.15
+ 0.5 2.16
+ 0.5 2.17
+ 0.5 2.18
+ 0.5 2.19
+ 0.5 2.2
+ 0.5 2.21
+ 0.5 2.22
+ 0.5 2.23
+ 0.5 2.24
+ 0.5 2.25
+ 0.5 2.26
+ 0.5 2.27
+ 0.5 2.28
+ 0.5 2.29
+ 0.5 2.3
+ 0.5 2.31
+ 0.5 2.32
+ 0.5 2.33
+ 0.5 2.34
+ 0.5 2.35
+ 0.5 2.36
+ 0.5 2.37
+ 0.5 2.38
+ 0.5 2.39
+ 0.5 2.4
+ 0.5 2.41
+ 0.5 2.42
+ 0.5 2.43
+ 0.5 2.44
+ 0.5 2.45
+ 0.5 2.46
+ 0.5 2.47
+ 0.5 2.48
+ 0.5 2.49
+ 0.5 2.5
+ 0.51 1.25
+ 0.51 1.26
+ 0.51 1.27
+ 0.51 1.28
+ 0.51 1.29
+ 0.51 1.3
+ 0.51 1.31
+ 0.51 1.32
+ 0.51 1.33
+ 0.51 1.34
+ 0.51 1.35
+ 0.51 1.36
+ 0.51 1.37
+ 0.51 1.38
+ 0.51 1.39
+ 0.51 1.4
+ 0.51 1.41
+ 0.51 1.42
+ 0.51 1.43
+ 0.51 1.44
+ 0.51 1.45
+ 0.51 1.46
+ 0.51 1.47
+ 0.51 1.48
+ 0.51 1.49
+ 0.51 1.5
+ 0.51 1.51
+ 0.51 1.52
+ 0.51 1.53
+ 0.51 1.54
+ 0.51 1.55
+ 0.51 1.56
+ 0.51 1.57
+ 0.51 1.58
+ 0.51 1.59
+ 0.51 1.6
+ 0.51 1.61
+ 0.51 1.62
+ 0.51 1.63
+ 0.51 1.64
+ 0.51 1.65
+ 0.51 1.66
+ 0.51 1.67
+ 0.51 1.68
+ 0.51 1.69
+ 0.51 1.7
+ 0.51 1.71
+ 0.51 1.72
+ 0.51 1.73
+ 0.51 1.74
+ 0.51 1.75
+ 0.51 1.76
+ 0.51 1.77
+ 0.51 1.78
+ 0.51 1.79
+ 0.51 1.8
+ 0.51 1.81
+ 0.51 1.82
+ 0.51 1.83
+ 0.51 1.84
+ 0.51 1.85
+ 0.51 1.86
+ 0.51 1.87
+ 0.51 1.88
+ 0.51 1.89
+ 0.51 1.9
+ 0.51 1.91
+ 0.51 1.92
+ 0.51 1.93
+ 0.51 1.94
+ 0.51 1.95
+ 0.51 1.96
+ 0.51 1.97
+ 0.51 1.98
+ 0.51 1.99
+ 0.51 2.0
+ 0.51 2.01
+ 0.51 2.02
+ 0.51 2.03
+ 0.51 2.04
+ 0.51 2.05
+ 0.51 2.06
+ 0.51 2.07
+ 0.51 2.08
+ 0.51 2.09
+ 0.51 2.1
+ 0.51 2.11
+ 0.51 2.12
+ 0.51 2.13
+ 0.51 2.14
+ 0.51 2.15
+ 0.51 2.16
+ 0.51 2.17
+ 0.51 2.18
+ 0.51 2.19
+ 0.51 2.2
+ 0.51 2.21
+ 0.51 2.22
+ 0.51 2.23
+ 0.51 2.24
+ 0.51 2.25
+ 0.51 2.26
+ 0.51 2.27
+ 0.51 2.28
+ 0.51 2.29
+ 0.51 2.3
+ 0.51 2.31
+ 0.51 2.32
+ 0.51 2.33
+ 0.51 2.34
+ 0.51 2.35
+ 0.51 2.36
+ 0.51 2.37
+ 0.51 2.38
+ 0.51 2.39
+ 0.51 2.4
+ 0.51 2.41
+ 0.51 2.42
+ 0.51 2.43
+ 0.51 2.44
+ 0.51 2.45
+ 0.51 2.46
+ 0.51 2.47
+ 0.51 2.48
+ 0.51 2.49
+ 0.51 2.5
+ 0.52 1.25
+ 0.52 1.26
+ 0.52 1.27
+ 0.52 1.28
+ 0.52 1.29
+ 0.52 1.3
+ 0.52 1.31
+ 0.52 1.32
+ 0.52 1.33
+ 0.52 1.34
+ 0.52 1.35
+ 0.52 1.36
+ 0.52 1.37
+ 0.52 1.38
+ 0.52 1.39
+ 0.52 1.4
+ 0.52 1.41
+ 0.52 1.42
+ 0.52 1.43
+ 0.52 1.44
+ 0.52 1.45
+ 0.52 1.46
+ 0.52 1.47
+ 0.52 1.48
+ 0.52 1.49
+ 0.52 1.5
+ 0.52 1.51
+ 0.52 1.52
+ 0.52 1.53
+ 0.52 1.54
+ 0.52 1.55
+ 0.52 1.56
+ 0.52 1.57
+ 0.52 1.58
+ 0.52 1.59
+ 0.52 1.6
+ 0.52 1.61
+ 0.52 1.62
+ 0.52 1.63
+ 0.52 1.64
+ 0.52 1.65
+ 0.52 1.66
+ 0.52 1.67
+ 0.52 1.68
+ 0.52 1.69
+ 0.52 1.7
+ 0.52 1.71
+ 0.52 1.72
+ 0.52 1.73
+ 0.52 1.74
+ 0.52 1.75
+ 0.52 1.76
+ 0.52 1.77
+ 0.52 1.78
+ 0.52 1.79
+ 0.52 1.8
+ 0.52 1.81
+ 0.52 1.82
+ 0.52 1.83
+ 0.52 1.84
+ 0.52 1.85
+ 0.52 1.86
+ 0.52 1.87
+ 0.52 1.88
+ 0.52 1.89
+ 0.52 1.9
+ 0.52 1.91
+ 0.52 1.92
+ 0.52 1.93
+ 0.52 1.94
+ 0.52 1.95
+ 0.52 1.96
+ 0.52 1.97
+ 0.52 1.98
+ 0.52 1.99
+ 0.52 2.0
+ 0.52 2.01
+ 0.52 2.02
+ 0.52 2.03
+ 0.52 2.04
+ 0.52 2.05
+ 0.52 2.06
+ 0.52 2.07
+ 0.52 2.08
+ 0.52 2.09
+ 0.52 2.1
+ 0.52 2.11
+ 0.52 2.12
+ 0.52 2.13
+ 0.52 2.14
+ 0.52 2.15
+ 0.52 2.16
+ 0.52 2.17
+ 0.52 2.18
+ 0.52 2.19
+ 0.52 2.2
+ 0.52 2.21
+ 0.52 2.22
+ 0.52 2.23
+ 0.52 2.24
+ 0.52 2.25
+ 0.52 2.26
+ 0.52 2.27
+ 0.52 2.28
+ 0.52 2.29
+ 0.52 2.3
+ 0.52 2.31
+ 0.52 2.32
+ 0.52 2.33
+ 0.52 2.34
+ 0.52 2.35
+ 0.52 2.36
+ 0.52 2.37
+ 0.52 2.38
+ 0.52 2.39
+ 0.52 2.4
+ 0.52 2.41
+ 0.52 2.42
+ 0.52 2.43
+ 0.52 2.44
+ 0.52 2.45
+ 0.52 2.46
+ 0.52 2.47
+ 0.52 2.48
+ 0.52 2.49
+ 0.52 2.5
+ 0.53 1.25
+ 0.53 1.26
+ 0.53 1.27
+ 0.53 1.28
+ 0.53 1.29
+ 0.53 1.3
+ 0.53 1.31
+ 0.53 1.32
+ 0.53 1.33
+ 0.53 1.34
+ 0.53 1.35
+ 0.53 1.36
+ 0.53 1.37
+ 0.53 1.38
+ 0.53 1.39
+ 0.53 1.4
+ 0.53 1.41
+ 0.53 1.42
+ 0.53 1.43
+ 0.53 1.44
+ 0.53 1.45
+ 0.53 1.46
+ 0.53 1.47
+ 0.53 1.48
+ 0.53 1.49
+ 0.53 1.5
+ 0.53 1.51
+ 0.53 1.52
+ 0.53 1.53
+ 0.53 1.54
+ 0.53 1.55
+ 0.53 1.56
+ 0.53 1.57
+ 0.53 1.58
+ 0.53 1.59
+ 0.53 1.6
+ 0.53 1.61
+ 0.53 1.62
+ 0.53 1.63
+ 0.53 1.64
+ 0.53 1.65
+ 0.53 1.66
+ 0.53 1.67
+ 0.53 1.68
+ 0.53 1.69
+ 0.53 1.7
+ 0.53 1.71
+ 0.53 1.72
+ 0.53 1.73
+ 0.53 1.74
+ 0.53 1.75
+ 0.53 1.76
+ 0.53 1.77
+ 0.53 1.78
+ 0.53 1.79
+ 0.53 1.8
+ 0.53 1.81
+ 0.53 1.82
+ 0.53 1.83
+ 0.53 1.84
+ 0.53 1.85
+ 0.53 1.86
+ 0.53 1.87
+ 0.53 1.88
+ 0.53 1.89
+ 0.53 1.9
+ 0.53 1.91
+ 0.53 1.92
+ 0.53 1.93
+ 0.53 1.94
+ 0.53 1.95
+ 0.53 1.96
+ 0.53 1.97
+ 0.53 1.98
+ 0.53 1.99
+ 0.53 2.0
+ 0.53 2.01
+ 0.53 2.02
+ 0.53 2.03
+ 0.53 2.04
+ 0.53 2.05
+ 0.53 2.06
+ 0.53 2.07
+ 0.53 2.08
+ 0.53 2.09
+ 0.53 2.1
+ 0.53 2.11
+ 0.53 2.12
+ 0.53 2.13
+ 0.53 2.14
+ 0.53 2.15
+ 0.53 2.16
+ 0.53 2.17
+ 0.53 2.18
+ 0.53 2.19
+ 0.53 2.2
+ 0.53 2.21
+ 0.53 2.22
+ 0.53 2.23
+ 0.53 2.24
+ 0.53 2.25
+ 0.53 2.26
+ 0.53 2.27
+ 0.53 2.28
+ 0.53 2.29
+ 0.53 2.3
+ 0.53 2.31
+ 0.53 2.32
+ 0.53 2.33
+ 0.53 2.34
+ 0.53 2.35
+ 0.53 2.36
+ 0.53 2.37
+ 0.53 2.38
+ 0.53 2.39
+ 0.53 2.4
+ 0.53 2.41
+ 0.53 2.42
+ 0.53 2.43
+ 0.53 2.44
+ 0.53 2.45
+ 0.53 2.46
+ 0.53 2.47
+ 0.53 2.48
+ 0.53 2.49
+ 0.53 2.5
+ 0.54 1.25
+ 0.54 1.26
+ 0.54 1.27
+ 0.54 1.28
+ 0.54 1.29
+ 0.54 1.3
+ 0.54 1.31
+ 0.54 1.32
+ 0.54 1.33
+ 0.54 1.34
+ 0.54 1.35
+ 0.54 1.36
+ 0.54 1.37
+ 0.54 1.38
+ 0.54 1.39
+ 0.54 1.4
+ 0.54 1.41
+ 0.54 1.42
+ 0.54 1.43
+ 0.54 1.44
+ 0.54 1.45
+ 0.54 1.46
+ 0.54 1.47
+ 0.54 1.48
+ 0.54 1.49
+ 0.54 1.5
+ 0.54 1.51
+ 0.54 1.52
+ 0.54 1.53
+ 0.54 1.54
+ 0.54 1.55
+ 0.54 1.56
+ 0.54 1.57
+ 0.54 1.58
+ 0.54 1.59
+ 0.54 1.6
+ 0.54 1.61
+ 0.54 1.62
+ 0.54 1.63
+ 0.54 1.64
+ 0.54 1.65
+ 0.54 1.66
+ 0.54 1.67
+ 0.54 1.68
+ 0.54 1.69
+ 0.54 1.7
+ 0.54 1.71
+ 0.54 1.72
+ 0.54 1.73
+ 0.54 1.74
+ 0.54 1.75
+ 0.54 1.76
+ 0.54 1.77
+ 0.54 1.78
+ 0.54 1.79
+ 0.54 1.8
+ 0.54 1.81
+ 0.54 1.82
+ 0.54 1.83
+ 0.54 1.84
+ 0.54 1.85
+ 0.54 1.86
+ 0.54 1.87
+ 0.54 1.88
+ 0.54 1.89
+ 0.54 1.9
+ 0.54 1.91
+ 0.54 1.92
+ 0.54 1.93
+ 0.54 1.94
+ 0.54 1.95
+ 0.54 1.96
+ 0.54 1.97
+ 0.54 1.98
+ 0.54 1.99
+ 0.54 2.0
+ 0.54 2.01
+ 0.54 2.02
+ 0.54 2.03
+ 0.54 2.04
+ 0.54 2.05
+ 0.54 2.06
+ 0.54 2.07
+ 0.54 2.08
+ 0.54 2.09
+ 0.54 2.1
+ 0.54 2.11
+ 0.54 2.12
+ 0.54 2.13
+ 0.54 2.14
+ 0.54 2.15
+ 0.54 2.16
+ 0.54 2.17
+ 0.54 2.18
+ 0.54 2.19
+ 0.54 2.2
+ 0.54 2.21
+ 0.54 2.22
+ 0.54 2.23
+ 0.54 2.24
+ 0.54 2.25
+ 0.54 2.26
+ 0.54 2.27
+ 0.54 2.28
+ 0.54 2.29
+ 0.54 2.3
+ 0.54 2.31
+ 0.54 2.32
+ 0.54 2.33
+ 0.54 2.34
+ 0.54 2.35
+ 0.54 2.36
+ 0.54 2.37
+ 0.54 2.38
+ 0.54 2.39
+ 0.54 2.4
+ 0.54 2.41
+ 0.54 2.42
+ 0.54 2.43
+ 0.54 2.44
+ 0.54 2.45
+ 0.54 2.46
+ 0.54 2.47
+ 0.54 2.48
+ 0.54 2.49
+ 0.54 2.5
+ 0.55 1.25
+ 0.55 1.26
+ 0.55 1.27
+ 0.55 1.28
+ 0.55 1.29
+ 0.55 1.3
+ 0.55 1.31
+ 0.55 1.32
+ 0.55 1.33
+ 0.55 1.34
+ 0.55 1.35
+ 0.55 1.36
+ 0.55 1.37
+ 0.55 1.38
+ 0.55 1.39
+ 0.55 1.4
+ 0.55 1.41
+ 0.55 1.42
+ 0.55 1.43
+ 0.55 1.44
+ 0.55 1.45
+ 0.55 1.46
+ 0.55 1.47
+ 0.55 1.48
+ 0.55 1.49
+ 0.55 1.5
+ 0.55 1.51
+ 0.55 1.52
+ 0.55 1.53
+ 0.55 1.54
+ 0.55 1.55
+ 0.55 1.56
+ 0.55 1.57
+ 0.55 1.58
+ 0.55 1.59
+ 0.55 1.6
+ 0.55 1.61
+ 0.55 1.62
+ 0.55 1.63
+ 0.55 1.64
+ 0.55 1.65
+ 0.55 1.66
+ 0.55 1.67
+ 0.55 1.68
+ 0.55 1.69
+ 0.55 1.7
+ 0.55 1.71
+ 0.55 1.72
+ 0.55 1.73
+ 0.55 1.74
+ 0.55 1.75
+ 0.55 1.76
+ 0.55 1.77
+ 0.55 1.78
+ 0.55 1.79
+ 0.55 1.8
+ 0.55 1.81
+ 0.55 1.82
+ 0.55 1.83
+ 0.55 1.84
+ 0.55 1.85
+ 0.55 1.86
+ 0.55 1.87
+ 0.55 1.88
+ 0.55 1.89
+ 0.55 1.9
+ 0.55 1.91
+ 0.55 1.92
+ 0.55 1.93
+ 0.55 1.94
+ 0.55 1.95
+ 0.55 1.96
+ 0.55 1.97
+ 0.55 1.98
+ 0.55 1.99
+ 0.55 2.0
+ 0.55 2.01
+ 0.55 2.02
+ 0.55 2.03
+ 0.55 2.04
+ 0.55 2.05
+ 0.55 2.06
+ 0.55 2.07
+ 0.55 2.08
+ 0.55 2.09
+ 0.55 2.1
+ 0.55 2.11
+ 0.55 2.12
+ 0.55 2.13
+ 0.55 2.14
+ 0.55 2.15
+ 0.55 2.16
+ 0.55 2.17
+ 0.55 2.18
+ 0.55 2.19
+ 0.55 2.2
+ 0.55 2.21
+ 0.55 2.22
+ 0.55 2.23
+ 0.55 2.24
+ 0.55 2.25
+ 0.55 2.26
+ 0.55 2.27
+ 0.55 2.28
+ 0.55 2.29
+ 0.55 2.3
+ 0.55 2.31
+ 0.55 2.32
+ 0.55 2.33
+ 0.55 2.34
+ 0.55 2.35
+ 0.55 2.36
+ 0.55 2.37
+ 0.55 2.38
+ 0.55 2.39
+ 0.55 2.4
+ 0.55 2.41
+ 0.55 2.42
+ 0.55 2.43
+ 0.55 2.44
+ 0.55 2.45
+ 0.55 2.46
+ 0.55 2.47
+ 0.55 2.48
+ 0.55 2.49
+ 0.55 2.5
+ 0.56 1.25
+ 0.56 1.26
+ 0.56 1.27
+ 0.56 1.28
+ 0.56 1.29
+ 0.56 1.3
+ 0.56 1.31
+ 0.56 1.32
+ 0.56 1.33
+ 0.56 1.34
+ 0.56 1.35
+ 0.56 1.36
+ 0.56 1.37
+ 0.56 1.38
+ 0.56 1.39
+ 0.56 1.4
+ 0.56 1.41
+ 0.56 1.42
+ 0.56 1.43
+ 0.56 1.44
+ 0.56 1.45
+ 0.56 1.46
+ 0.56 1.47
+ 0.56 1.48
+ 0.56 1.49
+ 0.56 1.5
+ 0.56 1.51
+ 0.56 1.52
+ 0.56 1.53
+ 0.56 1.54
+ 0.56 1.55
+ 0.56 1.56
+ 0.56 1.57
+ 0.56 1.58
+ 0.56 1.59
+ 0.56 1.6
+ 0.56 1.61
+ 0.56 1.62
+ 0.56 1.63
+ 0.56 1.64
+ 0.56 1.65
+ 0.56 1.66
+ 0.56 1.67
+ 0.56 1.68
+ 0.56 1.69
+ 0.56 1.7
+ 0.56 1.71
+ 0.56 1.72
+ 0.56 1.73
+ 0.56 1.74
+ 0.56 1.75
+ 0.56 1.76
+ 0.56 1.77
+ 0.56 1.78
+ 0.56 1.79
+ 0.56 1.8
+ 0.56 1.81
+ 0.56 1.82
+ 0.56 1.83
+ 0.56 1.84
+ 0.56 1.85
+ 0.56 1.86
+ 0.56 1.87
+ 0.56 1.88
+ 0.56 1.89
+ 0.56 1.9
+ 0.56 1.91
+ 0.56 1.92
+ 0.56 1.93
+ 0.56 1.94
+ 0.56 1.95
+ 0.56 1.96
+ 0.56 1.97
+ 0.56 1.98
+ 0.56 1.99
+ 0.56 2.0
+ 0.56 2.01
+ 0.56 2.02
+ 0.56 2.03
+ 0.56 2.04
+ 0.56 2.05
+ 0.56 2.06
+ 0.56 2.07
+ 0.56 2.08
+ 0.56 2.09
+ 0.56 2.1
+ 0.56 2.11
+ 0.56 2.12
+ 0.56 2.13
+ 0.56 2.14
+ 0.56 2.15
+ 0.56 2.16
+ 0.56 2.17
+ 0.56 2.18
+ 0.56 2.19
+ 0.56 2.2
+ 0.56 2.21
+ 0.56 2.22
+ 0.56 2.23
+ 0.56 2.24
+ 0.56 2.25
+ 0.56 2.26
+ 0.56 2.27
+ 0.56 2.28
+ 0.56 2.29
+ 0.56 2.3
+ 0.56 2.31
+ 0.56 2.32
+ 0.56 2.33
+ 0.56 2.34
+ 0.56 2.35
+ 0.56 2.36
+ 0.56 2.37
+ 0.56 2.38
+ 0.56 2.39
+ 0.56 2.4
+ 0.56 2.41
+ 0.56 2.42
+ 0.56 2.43
+ 0.56 2.44
+ 0.56 2.45
+ 0.56 2.46
+ 0.56 2.47
+ 0.56 2.48
+ 0.56 2.49
+ 0.56 2.5
+ 0.57 1.25
+ 0.57 1.26
+ 0.57 1.27
+ 0.57 1.28
+ 0.57 1.29
+ 0.57 1.3
+ 0.57 1.31
+ 0.57 1.32
+ 0.57 1.33
+ 0.57 1.34
+ 0.57 1.35
+ 0.57 1.36
+ 0.57 1.37
+ 0.57 1.38
+ 0.57 1.39
+ 0.57 1.4
+ 0.57 1.41
+ 0.57 1.42
+ 0.57 1.43
+ 0.57 1.44
+ 0.57 1.45
+ 0.57 1.46
+ 0.57 1.47
+ 0.57 1.48
+ 0.57 1.49
+ 0.57 1.5
+ 0.57 1.51
+ 0.57 1.52
+ 0.57 1.53
+ 0.57 1.54
+ 0.57 1.55
+ 0.57 1.56
+ 0.57 1.57
+ 0.57 1.58
+ 0.57 1.59
+ 0.57 1.6
+ 0.57 1.61
+ 0.57 1.62
+ 0.57 1.63
+ 0.57 1.64
+ 0.57 1.65
+ 0.57 1.66
+ 0.57 1.67
+ 0.57 1.68
+ 0.57 1.69
+ 0.57 1.7
+ 0.57 1.71
+ 0.57 1.72
+ 0.57 1.73
+ 0.57 1.74
+ 0.57 1.75
+ 0.57 1.76
+ 0.57 1.77
+ 0.57 1.78
+ 0.57 1.79
+ 0.57 1.8
+ 0.57 1.81
+ 0.57 1.82
+ 0.57 1.83
+ 0.57 1.84
+ 0.57 1.85
+ 0.57 1.86
+ 0.57 1.87
+ 0.57 1.88
+ 0.57 1.89
+ 0.57 1.9
+ 0.57 1.91
+ 0.57 1.92
+ 0.57 1.93
+ 0.57 1.94
+ 0.57 1.95
+ 0.57 1.96
+ 0.57 1.97
+ 0.57 1.98
+ 0.57 1.99
+ 0.57 2.0
+ 0.57 2.01
+ 0.57 2.02
+ 0.57 2.03
+ 0.57 2.04
+ 0.57 2.05
+ 0.57 2.06
+ 0.57 2.07
+ 0.57 2.08
+ 0.57 2.09
+ 0.57 2.1
+ 0.57 2.11
+ 0.57 2.12
+ 0.57 2.13
+ 0.57 2.14
+ 0.57 2.15
+ 0.57 2.16
+ 0.57 2.17
+ 0.57 2.18
+ 0.57 2.19
+ 0.57 2.2
+ 0.57 2.21
+ 0.57 2.22
+ 0.57 2.23
+ 0.57 2.24
+ 0.57 2.25
+ 0.57 2.26
+ 0.57 2.27
+ 0.57 2.28
+ 0.57 2.29
+ 0.57 2.3
+ 0.57 2.31
+ 0.57 2.32
+ 0.57 2.33
+ 0.57 2.34
+ 0.57 2.35
+ 0.57 2.36
+ 0.57 2.37
+ 0.57 2.38
+ 0.57 2.39
+ 0.57 2.4
+ 0.57 2.41
+ 0.57 2.42
+ 0.57 2.43
+ 0.57 2.44
+ 0.57 2.45
+ 0.57 2.46
+ 0.57 2.47
+ 0.57 2.48
+ 0.57 2.49
+ 0.57 2.5
+ 0.58 1.25
+ 0.58 1.26
+ 0.58 1.27
+ 0.58 1.28
+ 0.58 1.29
+ 0.58 1.3
+ 0.58 1.31
+ 0.58 1.32
+ 0.58 1.33
+ 0.58 1.34
+ 0.58 1.35
+ 0.58 1.36
+ 0.58 1.37
+ 0.58 1.38
+ 0.58 1.39
+ 0.58 1.4
+ 0.58 1.41
+ 0.58 1.42
+ 0.58 1.43
+ 0.58 1.44
+ 0.58 1.45
+ 0.58 1.46
+ 0.58 1.47
+ 0.58 1.48
+ 0.58 1.49
+ 0.58 1.5
+ 0.58 1.51
+ 0.58 1.52
+ 0.58 1.53
+ 0.58 1.54
+ 0.58 1.55
+ 0.58 1.56
+ 0.58 1.57
+ 0.58 1.58
+ 0.58 1.59
+ 0.58 1.6
+ 0.58 1.61
+ 0.58 1.62
+ 0.58 1.63
+ 0.58 1.64
+ 0.58 1.65
+ 0.58 1.66
+ 0.58 1.67
+ 0.58 1.68
+ 0.58 1.69
+ 0.58 1.7
+ 0.58 1.71
+ 0.58 1.72
+ 0.58 1.73
+ 0.58 1.74
+ 0.58 1.75
+ 0.58 1.76
+ 0.58 1.77
+ 0.58 1.78
+ 0.58 1.79
+ 0.58 1.8
+ 0.58 1.81
+ 0.58 1.82
+ 0.58 1.83
+ 0.58 1.84
+ 0.58 1.85
+ 0.58 1.86
+ 0.58 1.87
+ 0.58 1.88
+ 0.58 1.89
+ 0.58 1.9
+ 0.58 1.91
+ 0.58 1.92
+ 0.58 1.93
+ 0.58 1.94
+ 0.58 1.95
+ 0.58 1.96
+ 0.58 1.97
+ 0.58 1.98
+ 0.58 1.99
+ 0.58 2.0
+ 0.58 2.01
+ 0.58 2.02
+ 0.58 2.03
+ 0.58 2.04
+ 0.58 2.05
+ 0.58 2.06
+ 0.58 2.07
+ 0.58 2.08
+ 0.58 2.09
+ 0.58 2.1
+ 0.58 2.11
+ 0.58 2.12
+ 0.58 2.13
+ 0.58 2.14
+ 0.58 2.15
+ 0.58 2.16
+ 0.58 2.17
+ 0.58 2.18
+ 0.58 2.19
+ 0.58 2.2
+ 0.58 2.21
+ 0.58 2.22
+ 0.58 2.23
+ 0.58 2.24
+ 0.58 2.25
+ 0.58 2.26
+ 0.58 2.27
+ 0.58 2.28
+ 0.58 2.29
+ 0.58 2.3
+ 0.58 2.31
+ 0.58 2.32
+ 0.58 2.33
+ 0.58 2.34
+ 0.58 2.35
+ 0.58 2.36
+ 0.58 2.37
+ 0.58 2.38
+ 0.58 2.39
+ 0.58 2.4
+ 0.58 2.41
+ 0.58 2.42
+ 0.58 2.43
+ 0.58 2.44
+ 0.58 2.45
+ 0.58 2.46
+ 0.58 2.47
+ 0.58 2.48
+ 0.58 2.49
+ 0.58 2.5
+ 0.59 1.25
+ 0.59 1.26
+ 0.59 1.27
+ 0.59 1.28
+ 0.59 1.29
+ 0.59 1.3
+ 0.59 1.31
+ 0.59 1.32
+ 0.59 1.33
+ 0.59 1.34
+ 0.59 1.35
+ 0.59 1.36
+ 0.59 1.37
+ 0.59 1.38
+ 0.59 1.39
+ 0.59 1.4
+ 0.59 1.41
+ 0.59 1.42
+ 0.59 1.43
+ 0.59 1.44
+ 0.59 1.45
+ 0.59 1.46
+ 0.59 1.47
+ 0.59 1.48
+ 0.59 1.49
+ 0.59 1.5
+ 0.59 1.51
+ 0.59 1.52
+ 0.59 1.53
+ 0.59 1.54
+ 0.59 1.55
+ 0.59 1.56
+ 0.59 1.57
+ 0.59 1.58
+ 0.59 1.59
+ 0.59 1.6
+ 0.59 1.61
+ 0.59 1.62
+ 0.59 1.63
+ 0.59 1.64
+ 0.59 1.65
+ 0.59 1.66
+ 0.59 1.67
+ 0.59 1.68
+ 0.59 1.69
+ 0.59 1.7
+ 0.59 1.71
+ 0.59 1.72
+ 0.59 1.73
+ 0.59 1.74
+ 0.59 1.75
+ 0.59 1.76
+ 0.59 1.77
+ 0.59 1.78
+ 0.59 1.79
+ 0.59 1.8
+ 0.59 1.81
+ 0.59 1.82
+ 0.59 1.83
+ 0.59 1.84
+ 0.59 1.85
+ 0.59 1.86
+ 0.59 1.87
+ 0.59 1.88
+ 0.59 1.89
+ 0.59 1.9
+ 0.59 1.91
+ 0.59 1.92
+ 0.59 1.93
+ 0.59 1.94
+ 0.59 1.95
+ 0.59 1.96
+ 0.59 1.97
+ 0.59 1.98
+ 0.59 1.99
+ 0.59 2.0
+ 0.59 2.01
+ 0.59 2.02
+ 0.59 2.03
+ 0.59 2.04
+ 0.59 2.05
+ 0.59 2.06
+ 0.59 2.07
+ 0.59 2.08
+ 0.59 2.09
+ 0.59 2.1
+ 0.59 2.11
+ 0.59 2.12
+ 0.59 2.13
+ 0.59 2.14
+ 0.59 2.15
+ 0.59 2.16
+ 0.59 2.17
+ 0.59 2.18
+ 0.59 2.19
+ 0.59 2.2
+ 0.59 2.21
+ 0.59 2.22
+ 0.59 2.23
+ 0.59 2.24
+ 0.59 2.25
+ 0.59 2.26
+ 0.59 2.27
+ 0.59 2.28
+ 0.59 2.29
+ 0.59 2.3
+ 0.59 2.31
+ 0.59 2.32
+ 0.59 2.33
+ 0.59 2.34
+ 0.59 2.35
+ 0.59 2.36
+ 0.59 2.37
+ 0.59 2.38
+ 0.59 2.39
+ 0.59 2.4
+ 0.59 2.41
+ 0.59 2.42
+ 0.59 2.43
+ 0.59 2.44
+ 0.59 2.45
+ 0.59 2.46
+ 0.59 2.47
+ 0.59 2.48
+ 0.59 2.49
+ 0.59 2.5
+ 0.6 1.25
+ 0.6 1.26
+ 0.6 1.27
+ 0.6 1.28
+ 0.6 1.29
+ 0.6 1.3
+ 0.6 1.31
+ 0.6 1.32
+ 0.6 1.33
+ 0.6 1.34
+ 0.6 1.35
+ 0.6 1.36
+ 0.6 1.37
+ 0.6 1.38
+ 0.6 1.39
+ 0.6 1.4
+ 0.6 1.41
+ 0.6 1.42
+ 0.6 1.43
+ 0.6 1.44
+ 0.6 1.45
+ 0.6 1.46
+ 0.6 1.47
+ 0.6 1.48
+ 0.6 1.49
+ 0.6 1.5
+ 0.6 1.51
+ 0.6 1.52
+ 0.6 1.53
+ 0.6 1.54
+ 0.6 1.55
+ 0.6 1.56
+ 0.6 1.57
+ 0.6 1.58
+ 0.6 1.59
+ 0.6 1.6
+ 0.6 1.61
+ 0.6 1.62
+ 0.6 1.63
+ 0.6 1.64
+ 0.6 1.65
+ 0.6 1.66
+ 0.6 1.67
+ 0.6 1.68
+ 0.6 1.69
+ 0.6 1.7
+ 0.6 1.71
+ 0.6 1.72
+ 0.6 1.73
+ 0.6 1.74
+ 0.6 1.75
+ 0.6 1.76
+ 0.6 1.77
+ 0.6 1.78
+ 0.6 1.79
+ 0.6 1.8
+ 0.6 1.81
+ 0.6 1.82
+ 0.6 1.83
+ 0.6 1.84
+ 0.6 1.85
+ 0.6 1.86
+ 0.6 1.87
+ 0.6 1.88
+ 0.6 1.89
+ 0.6 1.9
+ 0.6 1.91
+ 0.6 1.92
+ 0.6 1.93
+ 0.6 1.94
+ 0.6 1.95
+ 0.6 1.96
+ 0.6 1.97
+ 0.6 1.98
+ 0.6 1.99
+ 0.6 2.0
+ 0.6 2.01
+ 0.6 2.02
+ 0.6 2.03
+ 0.6 2.04
+ 0.6 2.05
+ 0.6 2.06
+ 0.6 2.07
+ 0.6 2.08
+ 0.6 2.09
+ 0.6 2.1
+ 0.6 2.11
+ 0.6 2.12
+ 0.6 2.13
+ 0.6 2.14
+ 0.6 2.15
+ 0.6 2.16
+ 0.6 2.17
+ 0.6 2.18
+ 0.6 2.19
+ 0.6 2.2
+ 0.6 2.21
+ 0.6 2.22
+ 0.6 2.23
+ 0.6 2.24
+ 0.6 2.25
+ 0.6 2.26
+ 0.6 2.27
+ 0.6 2.28
+ 0.6 2.29
+ 0.6 2.3
+ 0.6 2.31
+ 0.6 2.32
+ 0.6 2.33
+ 0.6 2.34
+ 0.6 2.35
+ 0.6 2.36
+ 0.6 2.37
+ 0.6 2.38
+ 0.6 2.39
+ 0.6 2.4
+ 0.6 2.41
+ 0.6 2.42
+ 0.6 2.43
+ 0.6 2.44
+ 0.6 2.45
+ 0.6 2.46
+ 0.6 2.47
+ 0.6 2.48
+ 0.6 2.49
+ 0.6 2.5
+ 0.61 1.25
+ 0.61 1.26
+ 0.61 1.27
+ 0.61 1.28
+ 0.61 1.29
+ 0.61 1.3
+ 0.61 1.31
+ 0.61 1.32
+ 0.61 1.33
+ 0.61 1.34
+ 0.61 1.35
+ 0.61 1.36
+ 0.61 1.37
+ 0.61 1.38
+ 0.61 1.39
+ 0.61 1.4
+ 0.61 1.41
+ 0.61 1.42
+ 0.61 1.43
+ 0.61 1.44
+ 0.61 1.45
+ 0.61 1.46
+ 0.61 1.47
+ 0.61 1.48
+ 0.61 1.49
+ 0.61 1.5
+ 0.61 1.51
+ 0.61 1.52
+ 0.61 1.53
+ 0.61 1.54
+ 0.61 1.55
+ 0.61 1.56
+ 0.61 1.57
+ 0.61 1.58
+ 0.61 1.59
+ 0.61 1.6
+ 0.61 1.61
+ 0.61 1.62
+ 0.61 1.63
+ 0.61 1.64
+ 0.61 1.65
+ 0.61 1.66
+ 0.61 1.67
+ 0.61 1.68
+ 0.61 1.69
+ 0.61 1.7
+ 0.61 1.71
+ 0.61 1.72
+ 0.61 1.73
+ 0.61 1.74
+ 0.61 1.75
+ 0.61 1.76
+ 0.61 1.77
+ 0.61 1.78
+ 0.61 1.79
+ 0.61 1.8
+ 0.61 1.81
+ 0.61 1.82
+ 0.61 1.83
+ 0.61 1.84
+ 0.61 1.85
+ 0.61 1.86
+ 0.61 1.87
+ 0.61 1.88
+ 0.61 1.89
+ 0.61 1.9
+ 0.61 1.91
+ 0.61 1.92
+ 0.61 1.93
+ 0.61 1.94
+ 0.61 1.95
+ 0.61 1.96
+ 0.61 1.97
+ 0.61 1.98
+ 0.61 1.99
+ 0.61 2.0
+ 0.61 2.01
+ 0.61 2.02
+ 0.61 2.03
+ 0.61 2.04
+ 0.61 2.05
+ 0.61 2.06
+ 0.61 2.07
+ 0.61 2.08
+ 0.61 2.09
+ 0.61 2.1
+ 0.61 2.11
+ 0.61 2.12
+ 0.61 2.13
+ 0.61 2.14
+ 0.61 2.15
+ 0.61 2.16
+ 0.61 2.17
+ 0.61 2.18
+ 0.61 2.19
+ 0.61 2.2
+ 0.61 2.21
+ 0.61 2.22
+ 0.61 2.23
+ 0.61 2.24
+ 0.61 2.25
+ 0.61 2.26
+ 0.61 2.27
+ 0.61 2.28
+ 0.61 2.29
+ 0.61 2.3
+ 0.61 2.31
+ 0.61 2.32
+ 0.61 2.33
+ 0.61 2.34
+ 0.61 2.35
+ 0.61 2.36
+ 0.61 2.37
+ 0.61 2.38
+ 0.61 2.39
+ 0.61 2.4
+ 0.61 2.41
+ 0.61 2.42
+ 0.61 2.43
+ 0.61 2.44
+ 0.61 2.45
+ 0.61 2.46
+ 0.61 2.47
+ 0.61 2.48
+ 0.61 2.49
+ 0.61 2.5
+ 0.62 1.25
+ 0.62 1.26
+ 0.62 1.27
+ 0.62 1.28
+ 0.62 1.29
+ 0.62 1.3
+ 0.62 1.31
+ 0.62 1.32
+ 0.62 1.33
+ 0.62 1.34
+ 0.62 1.35
+ 0.62 1.36
+ 0.62 1.37
+ 0.62 1.38
+ 0.62 1.39
+ 0.62 1.4
+ 0.62 1.41
+ 0.62 1.42
+ 0.62 1.43
+ 0.62 1.44
+ 0.62 1.45
+ 0.62 1.46
+ 0.62 1.47
+ 0.62 1.48
+ 0.62 1.49
+ 0.62 1.5
+ 0.62 1.51
+ 0.62 1.52
+ 0.62 1.53
+ 0.62 1.54
+ 0.62 1.55
+ 0.62 1.56
+ 0.62 1.57
+ 0.62 1.58
+ 0.62 1.59
+ 0.62 1.6
+ 0.62 1.61
+ 0.62 1.62
+ 0.62 1.63
+ 0.62 1.64
+ 0.62 1.65
+ 0.62 1.66
+ 0.62 1.67
+ 0.62 1.68
+ 0.62 1.69
+ 0.62 1.7
+ 0.62 1.71
+ 0.62 1.72
+ 0.62 1.73
+ 0.62 1.74
+ 0.62 1.75
+ 0.62 1.76
+ 0.62 1.77
+ 0.62 1.78
+ 0.62 1.79
+ 0.62 1.8
+ 0.62 1.81
+ 0.62 1.82
+ 0.62 1.83
+ 0.62 1.84
+ 0.62 1.85
+ 0.62 1.86
+ 0.62 1.87
+ 0.62 1.88
+ 0.62 1.89
+ 0.62 1.9
+ 0.62 1.91
+ 0.62 1.92
+ 0.62 1.93
+ 0.62 1.94
+ 0.62 1.95
+ 0.62 1.96
+ 0.62 1.97
+ 0.62 1.98
+ 0.62 1.99
+ 0.62 2.0
+ 0.62 2.01
+ 0.62 2.02
+ 0.62 2.03
+ 0.62 2.04
+ 0.62 2.05
+ 0.62 2.06
+ 0.62 2.07
+ 0.62 2.08
+ 0.62 2.09
+ 0.62 2.1
+ 0.62 2.11
+ 0.62 2.12
+ 0.62 2.13
+ 0.62 2.14
+ 0.62 2.15
+ 0.62 2.16
+ 0.62 2.17
+ 0.62 2.18
+ 0.62 2.19
+ 0.62 2.2
+ 0.62 2.21
+ 0.62 2.22
+ 0.62 2.23
+ 0.62 2.24
+ 0.62 2.25
+ 0.62 2.26
+ 0.62 2.27
+ 0.62 2.28
+ 0.62 2.29
+ 0.62 2.3
+ 0.62 2.31
+ 0.62 2.32
+ 0.62 2.33
+ 0.62 2.34
+ 0.62 2.35
+ 0.62 2.36
+ 0.62 2.37
+ 0.62 2.38
+ 0.62 2.39
+ 0.62 2.4
+ 0.62 2.41
+ 0.62 2.42
+ 0.62 2.43
+ 0.62 2.44
+ 0.62 2.45
+ 0.62 2.46
+ 0.62 2.47
+ 0.62 2.48
+ 0.62 2.49
+ 0.62 2.5
+ 0.63 1.25
+ 0.63 1.26
+ 0.63 1.27
+ 0.63 1.28
+ 0.63 1.29
+ 0.63 1.3
+ 0.63 1.31
+ 0.63 1.32
+ 0.63 1.33
+ 0.63 1.34
+ 0.63 1.35
+ 0.63 1.36
+ 0.63 1.37
+ 0.63 1.38
+ 0.63 1.39
+ 0.63 1.4
+ 0.63 1.41
+ 0.63 1.42
+ 0.63 1.43
+ 0.63 1.44
+ 0.63 1.45
+ 0.63 1.46
+ 0.63 1.47
+ 0.63 1.48
+ 0.63 1.49
+ 0.63 1.5
+ 0.63 1.51
+ 0.63 1.52
+ 0.63 1.53
+ 0.63 1.54
+ 0.63 1.55
+ 0.63 1.56
+ 0.63 1.57
+ 0.63 1.58
+ 0.63 1.59
+ 0.63 1.6
+ 0.63 1.61
+ 0.63 1.62
+ 0.63 1.63
+ 0.63 1.64
+ 0.63 1.65
+ 0.63 1.66
+ 0.63 1.67
+ 0.63 1.68
+ 0.63 1.69
+ 0.63 1.7
+ 0.63 1.71
+ 0.63 1.72
+ 0.63 1.73
+ 0.63 1.74
+ 0.63 1.75
+ 0.63 1.76
+ 0.63 1.77
+ 0.63 1.78
+ 0.63 1.79
+ 0.63 1.8
+ 0.63 1.81
+ 0.63 1.82
+ 0.63 1.83
+ 0.63 1.84
+ 0.63 1.85
+ 0.63 1.86
+ 0.63 1.87
+ 0.63 1.88
+ 0.63 1.89
+ 0.63 1.9
+ 0.63 1.91
+ 0.63 1.92
+ 0.63 1.93
+ 0.63 1.94
+ 0.63 1.95
+ 0.63 1.96
+ 0.63 1.97
+ 0.63 1.98
+ 0.63 1.99
+ 0.63 2.0
+ 0.63 2.01
+ 0.63 2.02
+ 0.63 2.03
+ 0.63 2.04
+ 0.63 2.05
+ 0.63 2.06
+ 0.63 2.07
+ 0.63 2.08
+ 0.63 2.09
+ 0.63 2.1
+ 0.63 2.11
+ 0.63 2.12
+ 0.63 2.13
+ 0.63 2.14
+ 0.63 2.15
+ 0.63 2.16
+ 0.63 2.17
+ 0.63 2.18
+ 0.63 2.19
+ 0.63 2.2
+ 0.63 2.21
+ 0.63 2.22
+ 0.63 2.23
+ 0.63 2.24
+ 0.63 2.25
+ 0.63 2.26
+ 0.63 2.27
+ 0.63 2.28
+ 0.63 2.29
+ 0.63 2.3
+ 0.63 2.31
+ 0.63 2.32
+ 0.63 2.33
+ 0.63 2.34
+ 0.63 2.35
+ 0.63 2.36
+ 0.63 2.37
+ 0.63 2.38
+ 0.63 2.39
+ 0.63 2.4
+ 0.63 2.41
+ 0.63 2.42
+ 0.63 2.43
+ 0.63 2.44
+ 0.63 2.45
+ 0.63 2.46
+ 0.63 2.47
+ 0.63 2.48
+ 0.63 2.49
+ 0.63 2.5
+ 0.64 1.25
+ 0.64 1.26
+ 0.64 1.27
+ 0.64 1.28
+ 0.64 1.29
+ 0.64 1.3
+ 0.64 1.31
+ 0.64 1.32
+ 0.64 1.33
+ 0.64 1.34
+ 0.64 1.35
+ 0.64 1.36
+ 0.64 1.37
+ 0.64 1.38
+ 0.64 1.39
+ 0.64 1.4
+ 0.64 1.41
+ 0.64 1.42
+ 0.64 1.43
+ 0.64 1.44
+ 0.64 1.45
+ 0.64 1.46
+ 0.64 1.47
+ 0.64 1.48
+ 0.64 1.49
+ 0.64 1.5
+ 0.64 1.51
+ 0.64 1.52
+ 0.64 1.53
+ 0.64 1.54
+ 0.64 1.55
+ 0.64 1.56
+ 0.64 1.57
+ 0.64 1.58
+ 0.64 1.59
+ 0.64 1.6
+ 0.64 1.61
+ 0.64 1.62
+ 0.64 1.63
+ 0.64 1.64
+ 0.64 1.65
+ 0.64 1.66
+ 0.64 1.67
+ 0.64 1.68
+ 0.64 1.69
+ 0.64 1.7
+ 0.64 1.71
+ 0.64 1.72
+ 0.64 1.73
+ 0.64 1.74
+ 0.64 1.75
+ 0.64 1.76
+ 0.64 1.77
+ 0.64 1.78
+ 0.64 1.79
+ 0.64 1.8
+ 0.64 1.81
+ 0.64 1.82
+ 0.64 1.83
+ 0.64 1.84
+ 0.64 1.85
+ 0.64 1.86
+ 0.64 1.87
+ 0.64 1.88
+ 0.64 1.89
+ 0.64 1.9
+ 0.64 1.91
+ 0.64 1.92
+ 0.64 1.93
+ 0.64 1.94
+ 0.64 1.95
+ 0.64 1.96
+ 0.64 1.97
+ 0.64 1.98
+ 0.64 1.99
+ 0.64 2.0
+ 0.64 2.01
+ 0.64 2.02
+ 0.64 2.03
+ 0.64 2.04
+ 0.64 2.05
+ 0.64 2.06
+ 0.64 2.07
+ 0.64 2.08
+ 0.64 2.09
+ 0.64 2.1
+ 0.64 2.11
+ 0.64 2.12
+ 0.64 2.13
+ 0.64 2.14
+ 0.64 2.15
+ 0.64 2.16
+ 0.64 2.17
+ 0.64 2.18
+ 0.64 2.19
+ 0.64 2.2
+ 0.64 2.21
+ 0.64 2.22
+ 0.64 2.23
+ 0.64 2.24
+ 0.64 2.25
+ 0.64 2.26
+ 0.64 2.27
+ 0.64 2.28
+ 0.64 2.29
+ 0.64 2.3
+ 0.64 2.31
+ 0.64 2.32
+ 0.64 2.33
+ 0.64 2.34
+ 0.64 2.35
+ 0.64 2.36
+ 0.64 2.37
+ 0.64 2.38
+ 0.64 2.39
+ 0.64 2.4
+ 0.64 2.41
+ 0.64 2.42
+ 0.64 2.43
+ 0.64 2.44
+ 0.64 2.45
+ 0.64 2.46
+ 0.64 2.47
+ 0.64 2.48
+ 0.64 2.49
+ 0.64 2.5
+ 0.65 1.25
+ 0.65 1.26
+ 0.65 1.27
+ 0.65 1.28
+ 0.65 1.29
+ 0.65 1.3
+ 0.65 1.31
+ 0.65 1.32
+ 0.65 1.33
+ 0.65 1.34
+ 0.65 1.35
+ 0.65 1.36
+ 0.65 1.37
+ 0.65 1.38
+ 0.65 1.39
+ 0.65 1.4
+ 0.65 1.41
+ 0.65 1.42
+ 0.65 1.43
+ 0.65 1.44
+ 0.65 1.45
+ 0.65 1.46
+ 0.65 1.47
+ 0.65 1.48
+ 0.65 1.49
+ 0.65 1.5
+ 0.65 1.51
+ 0.65 1.52
+ 0.65 1.53
+ 0.65 1.54
+ 0.65 1.55
+ 0.65 1.56
+ 0.65 1.57
+ 0.65 1.58
+ 0.65 1.59
+ 0.65 1.6
+ 0.65 1.61
+ 0.65 1.62
+ 0.65 1.63
+ 0.65 1.64
+ 0.65 1.65
+ 0.65 1.66
+ 0.65 1.67
+ 0.65 1.68
+ 0.65 1.69
+ 0.65 1.7
+ 0.65 1.71
+ 0.65 1.72
+ 0.65 1.73
+ 0.65 1.74
+ 0.65 1.75
+ 0.65 1.76
+ 0.65 1.77
+ 0.65 1.78
+ 0.65 1.79
+ 0.65 1.8
+ 0.65 1.81
+ 0.65 1.82
+ 0.65 1.83
+ 0.65 1.84
+ 0.65 1.85
+ 0.65 1.86
+ 0.65 1.87
+ 0.65 1.88
+ 0.65 1.89
+ 0.65 1.9
+ 0.65 1.91
+ 0.65 1.92
+ 0.65 1.93
+ 0.65 1.94
+ 0.65 1.95
+ 0.65 1.96
+ 0.65 1.97
+ 0.65 1.98
+ 0.65 1.99
+ 0.65 2.0
+ 0.65 2.01
+ 0.65 2.02
+ 0.65 2.03
+ 0.65 2.04
+ 0.65 2.05
+ 0.65 2.06
+ 0.65 2.07
+ 0.65 2.08
+ 0.65 2.09
+ 0.65 2.1
+ 0.65 2.11
+ 0.65 2.12
+ 0.65 2.13
+ 0.65 2.14
+ 0.65 2.15
+ 0.65 2.16
+ 0.65 2.17
+ 0.65 2.18
+ 0.65 2.19
+ 0.65 2.2
+ 0.65 2.21
+ 0.65 2.22
+ 0.65 2.23
+ 0.65 2.24
+ 0.65 2.25
+ 0.65 2.26
+ 0.65 2.27
+ 0.65 2.28
+ 0.65 2.29
+ 0.65 2.3
+ 0.65 2.31
+ 0.65 2.32
+ 0.65 2.33
+ 0.65 2.34
+ 0.65 2.35
+ 0.65 2.36
+ 0.65 2.37
+ 0.65 2.38
+ 0.65 2.39
+ 0.65 2.4
+ 0.65 2.41
+ 0.65 2.42
+ 0.65 2.43
+ 0.65 2.44
+ 0.65 2.45
+ 0.65 2.46
+ 0.65 2.47
+ 0.65 2.48
+ 0.65 2.49
+ 0.65 2.5
+ 0.66 1.25
+ 0.66 1.26
+ 0.66 1.27
+ 0.66 1.28
+ 0.66 1.29
+ 0.66 1.3
+ 0.66 1.31
+ 0.66 1.32
+ 0.66 1.33
+ 0.66 1.34
+ 0.66 1.35
+ 0.66 1.36
+ 0.66 1.37
+ 0.66 1.38
+ 0.66 1.39
+ 0.66 1.4
+ 0.66 1.41
+ 0.66 1.42
+ 0.66 1.43
+ 0.66 1.44
+ 0.66 1.45
+ 0.66 1.46
+ 0.66 1.47
+ 0.66 1.48
+ 0.66 1.49
+ 0.66 1.5
+ 0.66 1.51
+ 0.66 1.52
+ 0.66 1.53
+ 0.66 1.54
+ 0.66 1.55
+ 0.66 1.56
+ 0.66 1.57
+ 0.66 1.58
+ 0.66 1.59
+ 0.66 1.6
+ 0.66 1.61
+ 0.66 1.62
+ 0.66 1.63
+ 0.66 1.64
+ 0.66 1.65
+ 0.66 1.66
+ 0.66 1.67
+ 0.66 1.68
+ 0.66 1.69
+ 0.66 1.7
+ 0.66 1.71
+ 0.66 1.72
+ 0.66 1.73
+ 0.66 1.74
+ 0.66 1.75
+ 0.66 1.76
+ 0.66 1.77
+ 0.66 1.78
+ 0.66 1.79
+ 0.66 1.8
+ 0.66 1.81
+ 0.66 1.82
+ 0.66 1.83
+ 0.66 1.84
+ 0.66 1.85
+ 0.66 1.86
+ 0.66 1.87
+ 0.66 1.88
+ 0.66 1.89
+ 0.66 1.9
+ 0.66 1.91
+ 0.66 1.92
+ 0.66 1.93
+ 0.66 1.94
+ 0.66 1.95
+ 0.66 1.96
+ 0.66 1.97
+ 0.66 1.98
+ 0.66 1.99
+ 0.66 2.0
+ 0.66 2.01
+ 0.66 2.02
+ 0.66 2.03
+ 0.66 2.04
+ 0.66 2.05
+ 0.66 2.06
+ 0.66 2.07
+ 0.66 2.08
+ 0.66 2.09
+ 0.66 2.1
+ 0.66 2.11
+ 0.66 2.12
+ 0.66 2.13
+ 0.66 2.14
+ 0.66 2.15
+ 0.66 2.16
+ 0.66 2.17
+ 0.66 2.18
+ 0.66 2.19
+ 0.66 2.2
+ 0.66 2.21
+ 0.66 2.22
+ 0.66 2.23
+ 0.66 2.24
+ 0.66 2.25
+ 0.66 2.26
+ 0.66 2.27
+ 0.66 2.28
+ 0.66 2.29
+ 0.66 2.3
+ 0.66 2.31
+ 0.66 2.32
+ 0.66 2.33
+ 0.66 2.34
+ 0.66 2.35
+ 0.66 2.36
+ 0.66 2.37
+ 0.66 2.38
+ 0.66 2.39
+ 0.66 2.4
+ 0.66 2.41
+ 0.66 2.42
+ 0.66 2.43
+ 0.66 2.44
+ 0.66 2.45
+ 0.66 2.46
+ 0.66 2.47
+ 0.66 2.48
+ 0.66 2.49
+ 0.66 2.5
+ 0.67 1.25
+ 0.67 1.26
+ 0.67 1.27
+ 0.67 1.28
+ 0.67 1.29
+ 0.67 1.3
+ 0.67 1.31
+ 0.67 1.32
+ 0.67 1.33
+ 0.67 1.34
+ 0.67 1.35
+ 0.67 1.36
+ 0.67 1.37
+ 0.67 1.38
+ 0.67 1.39
+ 0.67 1.4
+ 0.67 1.41
+ 0.67 1.42
+ 0.67 1.43
+ 0.67 1.44
+ 0.67 1.45
+ 0.67 1.46
+ 0.67 1.47
+ 0.67 1.48
+ 0.67 1.49
+ 0.67 1.5
+ 0.67 1.51
+ 0.67 1.52
+ 0.67 1.53
+ 0.67 1.54
+ 0.67 1.55
+ 0.67 1.56
+ 0.67 1.57
+ 0.67 1.58
+ 0.67 1.59
+ 0.67 1.6
+ 0.67 1.61
+ 0.67 1.62
+ 0.67 1.63
+ 0.67 1.64
+ 0.67 1.65
+ 0.67 1.66
+ 0.67 1.67
+ 0.67 1.68
+ 0.67 1.69
+ 0.67 1.7
+ 0.67 1.71
+ 0.67 1.72
+ 0.67 1.73
+ 0.67 1.74
+ 0.67 1.75
+ 0.67 1.76
+ 0.67 1.77
+ 0.67 1.78
+ 0.67 1.79
+ 0.67 1.8
+ 0.67 1.81
+ 0.67 1.82
+ 0.67 1.83
+ 0.67 1.84
+ 0.67 1.85
+ 0.67 1.86
+ 0.67 1.87
+ 0.67 1.88
+ 0.67 1.89
+ 0.67 1.9
+ 0.67 1.91
+ 0.67 1.92
+ 0.67 1.93
+ 0.67 1.94
+ 0.67 1.95
+ 0.67 1.96
+ 0.67 1.97
+ 0.67 1.98
+ 0.67 1.99
+ 0.67 2.0
+ 0.67 2.01
+ 0.67 2.02
+ 0.67 2.03
+ 0.67 2.04
+ 0.67 2.05
+ 0.67 2.06
+ 0.67 2.07
+ 0.67 2.08
+ 0.67 2.09
+ 0.67 2.1
+ 0.67 2.11
+ 0.67 2.12
+ 0.67 2.13
+ 0.67 2.14
+ 0.67 2.15
+ 0.67 2.16
+ 0.67 2.17
+ 0.67 2.18
+ 0.67 2.19
+ 0.67 2.2
+ 0.67 2.21
+ 0.67 2.22
+ 0.67 2.23
+ 0.67 2.24
+ 0.67 2.25
+ 0.67 2.26
+ 0.67 2.27
+ 0.67 2.28
+ 0.67 2.29
+ 0.67 2.3
+ 0.67 2.31
+ 0.67 2.32
+ 0.67 2.33
+ 0.67 2.34
+ 0.67 2.35
+ 0.67 2.36
+ 0.67 2.37
+ 0.67 2.38
+ 0.67 2.39
+ 0.67 2.4
+ 0.67 2.41
+ 0.67 2.42
+ 0.67 2.43
+ 0.67 2.44
+ 0.67 2.45
+ 0.67 2.46
+ 0.67 2.47
+ 0.67 2.48
+ 0.67 2.49
+ 0.67 2.5
+ 0.68 1.25
+ 0.68 1.26
+ 0.68 1.27
+ 0.68 1.28
+ 0.68 1.29
+ 0.68 1.3
+ 0.68 1.31
+ 0.68 1.32
+ 0.68 1.33
+ 0.68 1.34
+ 0.68 1.35
+ 0.68 1.36
+ 0.68 1.37
+ 0.68 1.38
+ 0.68 1.39
+ 0.68 1.4
+ 0.68 1.41
+ 0.68 1.42
+ 0.68 1.43
+ 0.68 1.44
+ 0.68 1.45
+ 0.68 1.46
+ 0.68 1.47
+ 0.68 1.48
+ 0.68 1.49
+ 0.68 1.5
+ 0.68 1.51
+ 0.68 1.52
+ 0.68 1.53
+ 0.68 1.54
+ 0.68 1.55
+ 0.68 1.56
+ 0.68 1.57
+ 0.68 1.58
+ 0.68 1.59
+ 0.68 1.6
+ 0.68 1.61
+ 0.68 1.62
+ 0.68 1.63
+ 0.68 1.64
+ 0.68 1.65
+ 0.68 1.66
+ 0.68 1.67
+ 0.68 1.68
+ 0.68 1.69
+ 0.68 1.7
+ 0.68 1.71
+ 0.68 1.72
+ 0.68 1.73
+ 0.68 1.74
+ 0.68 1.75
+ 0.68 1.76
+ 0.68 1.77
+ 0.68 1.78
+ 0.68 1.79
+ 0.68 1.8
+ 0.68 1.81
+ 0.68 1.82
+ 0.68 1.83
+ 0.68 1.84
+ 0.68 1.85
+ 0.68 1.86
+ 0.68 1.87
+ 0.68 1.88
+ 0.68 1.89
+ 0.68 1.9
+ 0.68 1.91
+ 0.68 1.92
+ 0.68 1.93
+ 0.68 1.94
+ 0.68 1.95
+ 0.68 1.96
+ 0.68 1.97
+ 0.68 1.98
+ 0.68 1.99
+ 0.68 2.0
+ 0.68 2.01
+ 0.68 2.02
+ 0.68 2.03
+ 0.68 2.04
+ 0.68 2.05
+ 0.68 2.06
+ 0.68 2.07
+ 0.68 2.08
+ 0.68 2.09
+ 0.68 2.1
+ 0.68 2.11
+ 0.68 2.12
+ 0.68 2.13
+ 0.68 2.14
+ 0.68 2.15
+ 0.68 2.16
+ 0.68 2.17
+ 0.68 2.18
+ 0.68 2.19
+ 0.68 2.2
+ 0.68 2.21
+ 0.68 2.22
+ 0.68 2.23
+ 0.68 2.24
+ 0.68 2.25
+ 0.68 2.26
+ 0.68 2.27
+ 0.68 2.28
+ 0.68 2.29
+ 0.68 2.3
+ 0.68 2.31
+ 0.68 2.32
+ 0.68 2.33
+ 0.68 2.34
+ 0.68 2.35
+ 0.68 2.36
+ 0.68 2.37
+ 0.68 2.38
+ 0.68 2.39
+ 0.68 2.4
+ 0.68 2.41
+ 0.68 2.42
+ 0.68 2.43
+ 0.68 2.44
+ 0.68 2.45
+ 0.68 2.46
+ 0.68 2.47
+ 0.68 2.48
+ 0.68 2.49
+ 0.68 2.5
+ 0.69 1.25
+ 0.69 1.26
+ 0.69 1.27
+ 0.69 1.28
+ 0.69 1.29
+ 0.69 1.3
+ 0.69 1.31
+ 0.69 1.32
+ 0.69 1.33
+ 0.69 1.34
+ 0.69 1.35
+ 0.69 1.36
+ 0.69 1.37
+ 0.69 1.38
+ 0.69 1.39
+ 0.69 1.4
+ 0.69 1.41
+ 0.69 1.42
+ 0.69 1.43
+ 0.69 1.44
+ 0.69 1.45
+ 0.69 1.46
+ 0.69 1.47
+ 0.69 1.48
+ 0.69 1.49
+ 0.69 1.5
+ 0.69 1.51
+ 0.69 1.52
+ 0.69 1.53
+ 0.69 1.54
+ 0.69 1.55
+ 0.69 1.56
+ 0.69 1.57
+ 0.69 1.58
+ 0.69 1.59
+ 0.69 1.6
+ 0.69 1.61
+ 0.69 1.62
+ 0.69 1.63
+ 0.69 1.64
+ 0.69 1.65
+ 0.69 1.66
+ 0.69 1.67
+ 0.69 1.68
+ 0.69 1.69
+ 0.69 1.7
+ 0.69 1.71
+ 0.69 1.72
+ 0.69 1.73
+ 0.69 1.74
+ 0.69 1.75
+ 0.69 1.76
+ 0.69 1.77
+ 0.69 1.78
+ 0.69 1.79
+ 0.69 1.8
+ 0.69 1.81
+ 0.69 1.82
+ 0.69 1.83
+ 0.69 1.84
+ 0.69 1.85
+ 0.69 1.86
+ 0.69 1.87
+ 0.69 1.88
+ 0.69 1.89
+ 0.69 1.9
+ 0.69 1.91
+ 0.69 1.92
+ 0.69 1.93
+ 0.69 1.94
+ 0.69 1.95
+ 0.69 1.96
+ 0.69 1.97
+ 0.69 1.98
+ 0.69 1.99
+ 0.69 2.0
+ 0.69 2.01
+ 0.69 2.02
+ 0.69 2.03
+ 0.69 2.04
+ 0.69 2.05
+ 0.69 2.06
+ 0.69 2.07
+ 0.69 2.08
+ 0.69 2.09
+ 0.69 2.1
+ 0.69 2.11
+ 0.69 2.12
+ 0.69 2.13
+ 0.69 2.14
+ 0.69 2.15
+ 0.69 2.16
+ 0.69 2.17
+ 0.69 2.18
+ 0.69 2.19
+ 0.69 2.2
+ 0.69 2.21
+ 0.69 2.22
+ 0.69 2.23
+ 0.69 2.24
+ 0.69 2.25
+ 0.69 2.26
+ 0.69 2.27
+ 0.69 2.28
+ 0.69 2.29
+ 0.69 2.3
+ 0.69 2.31
+ 0.69 2.32
+ 0.69 2.33
+ 0.69 2.34
+ 0.69 2.35
+ 0.69 2.36
+ 0.69 2.37
+ 0.69 2.38
+ 0.69 2.39
+ 0.69 2.4
+ 0.69 2.41
+ 0.69 2.42
+ 0.69 2.43
+ 0.69 2.44
+ 0.69 2.45
+ 0.69 2.46
+ 0.69 2.47
+ 0.69 2.48
+ 0.69 2.49
+ 0.69 2.5
+ 0.7 1.25
+ 0.7 1.26
+ 0.7 1.27
+ 0.7 1.28
+ 0.7 1.29
+ 0.7 1.3
+ 0.7 1.31
+ 0.7 1.32
+ 0.7 1.33
+ 0.7 1.34
+ 0.7 1.35
+ 0.7 1.36
+ 0.7 1.37
+ 0.7 1.38
+ 0.7 1.39
+ 0.7 1.4
+ 0.7 1.41
+ 0.7 1.42
+ 0.7 1.43
+ 0.7 1.44
+ 0.7 1.45
+ 0.7 1.46
+ 0.7 1.47
+ 0.7 1.48
+ 0.7 1.49
+ 0.7 1.5
+ 0.7 1.51
+ 0.7 1.52
+ 0.7 1.53
+ 0.7 1.54
+ 0.7 1.55
+ 0.7 1.56
+ 0.7 1.57
+ 0.7 1.58
+ 0.7 1.59
+ 0.7 1.6
+ 0.7 1.61
+ 0.7 1.62
+ 0.7 1.63
+ 0.7 1.64
+ 0.7 1.65
+ 0.7 1.66
+ 0.7 1.67
+ 0.7 1.68
+ 0.7 1.69
+ 0.7 1.7
+ 0.7 1.71
+ 0.7 1.72
+ 0.7 1.73
+ 0.7 1.74
+ 0.7 1.75
+ 0.7 1.76
+ 0.7 1.77
+ 0.7 1.78
+ 0.7 1.79
+ 0.7 1.8
+ 0.7 1.81
+ 0.7 1.82
+ 0.7 1.83
+ 0.7 1.84
+ 0.7 1.85
+ 0.7 1.86
+ 0.7 1.87
+ 0.7 1.88
+ 0.7 1.89
+ 0.7 1.9
+ 0.7 1.91
+ 0.7 1.92
+ 0.7 1.93
+ 0.7 1.94
+ 0.7 1.95
+ 0.7 1.96
+ 0.7 1.97
+ 0.7 1.98
+ 0.7 1.99
+ 0.7 2.0
+ 0.7 2.01
+ 0.7 2.02
+ 0.7 2.03
+ 0.7 2.04
+ 0.7 2.05
+ 0.7 2.06
+ 0.7 2.07
+ 0.7 2.08
+ 0.7 2.09
+ 0.7 2.1
+ 0.7 2.11
+ 0.7 2.12
+ 0.7 2.13
+ 0.7 2.14
+ 0.7 2.15
+ 0.7 2.16
+ 0.7 2.17
+ 0.7 2.18
+ 0.7 2.19
+ 0.7 2.2
+ 0.7 2.21
+ 0.7 2.22
+ 0.7 2.23
+ 0.7 2.24
+ 0.7 2.25
+ 0.7 2.26
+ 0.7 2.27
+ 0.7 2.28
+ 0.7 2.29
+ 0.7 2.3
+ 0.7 2.31
+ 0.7 2.32
+ 0.7 2.33
+ 0.7 2.34
+ 0.7 2.35
+ 0.7 2.36
+ 0.7 2.37
+ 0.7 2.38
+ 0.7 2.39
+ 0.7 2.4
+ 0.7 2.41
+ 0.7 2.42
+ 0.7 2.43
+ 0.7 2.44
+ 0.7 2.45
+ 0.7 2.46
+ 0.7 2.47
+ 0.7 2.48
+ 0.7 2.49
+ 0.7 2.5
+ 0.71 1.25
+ 0.71 1.26
+ 0.71 1.27
+ 0.71 1.28
+ 0.71 1.29
+ 0.71 1.3
+ 0.71 1.31
+ 0.71 1.32
+ 0.71 1.33
+ 0.71 1.34
+ 0.71 1.35
+ 0.71 1.36
+ 0.71 1.37
+ 0.71 1.38
+ 0.71 1.39
+ 0.71 1.4
+ 0.71 1.41
+ 0.71 1.42
+ 0.71 1.43
+ 0.71 1.44
+ 0.71 1.45
+ 0.71 1.46
+ 0.71 1.47
+ 0.71 1.48
+ 0.71 1.49
+ 0.71 1.5
+ 0.71 1.51
+ 0.71 1.52
+ 0.71 1.53
+ 0.71 1.54
+ 0.71 1.55
+ 0.71 1.56
+ 0.71 1.57
+ 0.71 1.58
+ 0.71 1.59
+ 0.71 1.6
+ 0.71 1.61
+ 0.71 1.62
+ 0.71 1.63
+ 0.71 1.64
+ 0.71 1.65
+ 0.71 1.66
+ 0.71 1.67
+ 0.71 1.68
+ 0.71 1.69
+ 0.71 1.7
+ 0.71 1.71
+ 0.71 1.72
+ 0.71 1.73
+ 0.71 1.74
+ 0.71 1.75
+ 0.71 1.76
+ 0.71 1.77
+ 0.71 1.78
+ 0.71 1.79
+ 0.71 1.8
+ 0.71 1.81
+ 0.71 1.82
+ 0.71 1.83
+ 0.71 1.84
+ 0.71 1.85
+ 0.71 1.86
+ 0.71 1.87
+ 0.71 1.88
+ 0.71 1.89
+ 0.71 1.9
+ 0.71 1.91
+ 0.71 1.92
+ 0.71 1.93
+ 0.71 1.94
+ 0.71 1.95
+ 0.71 1.96
+ 0.71 1.97
+ 0.71 1.98
+ 0.71 1.99
+ 0.71 2.0
+ 0.71 2.01
+ 0.71 2.02
+ 0.71 2.03
+ 0.71 2.04
+ 0.71 2.05
+ 0.71 2.06
+ 0.71 2.07
+ 0.71 2.08
+ 0.71 2.09
+ 0.71 2.1
+ 0.71 2.11
+ 0.71 2.12
+ 0.71 2.13
+ 0.71 2.14
+ 0.71 2.15
+ 0.71 2.16
+ 0.71 2.17
+ 0.71 2.18
+ 0.71 2.19
+ 0.71 2.2
+ 0.71 2.21
+ 0.71 2.22
+ 0.71 2.23
+ 0.71 2.24
+ 0.71 2.25
+ 0.71 2.26
+ 0.71 2.27
+ 0.71 2.28
+ 0.71 2.29
+ 0.71 2.3
+ 0.71 2.31
+ 0.71 2.32
+ 0.71 2.33
+ 0.71 2.34
+ 0.71 2.35
+ 0.71 2.36
+ 0.71 2.37
+ 0.71 2.38
+ 0.71 2.39
+ 0.71 2.4
+ 0.71 2.41
+ 0.71 2.42
+ 0.71 2.43
+ 0.71 2.44
+ 0.71 2.45
+ 0.71 2.46
+ 0.71 2.47
+ 0.71 2.48
+ 0.71 2.49
+ 0.71 2.5
+ 0.72 1.25
+ 0.72 1.26
+ 0.72 1.27
+ 0.72 1.28
+ 0.72 1.29
+ 0.72 1.3
+ 0.72 1.31
+ 0.72 1.32
+ 0.72 1.33
+ 0.72 1.34
+ 0.72 1.35
+ 0.72 1.36
+ 0.72 1.37
+ 0.72 1.38
+ 0.72 1.39
+ 0.72 1.4
+ 0.72 1.41
+ 0.72 1.42
+ 0.72 1.43
+ 0.72 1.44
+ 0.72 1.45
+ 0.72 1.46
+ 0.72 1.47
+ 0.72 1.48
+ 0.72 1.49
+ 0.72 1.5
+ 0.72 1.51
+ 0.72 1.52
+ 0.72 1.53
+ 0.72 1.54
+ 0.72 1.55
+ 0.72 1.56
+ 0.72 1.57
+ 0.72 1.58
+ 0.72 1.59
+ 0.72 1.6
+ 0.72 1.61
+ 0.72 1.62
+ 0.72 1.63
+ 0.72 1.64
+ 0.72 1.65
+ 0.72 1.66
+ 0.72 1.67
+ 0.72 1.68
+ 0.72 1.69
+ 0.72 1.7
+ 0.72 1.71
+ 0.72 1.72
+ 0.72 1.73
+ 0.72 1.74
+ 0.72 1.75
+ 0.72 1.76
+ 0.72 1.77
+ 0.72 1.78
+ 0.72 1.79
+ 0.72 1.8
+ 0.72 1.81
+ 0.72 1.82
+ 0.72 1.83
+ 0.72 1.84
+ 0.72 1.85
+ 0.72 1.86
+ 0.72 1.87
+ 0.72 1.88
+ 0.72 1.89
+ 0.72 1.9
+ 0.72 1.91
+ 0.72 1.92
+ 0.72 1.93
+ 0.72 1.94
+ 0.72 1.95
+ 0.72 1.96
+ 0.72 1.97
+ 0.72 1.98
+ 0.72 1.99
+ 0.72 2.0
+ 0.72 2.01
+ 0.72 2.02
+ 0.72 2.03
+ 0.72 2.04
+ 0.72 2.05
+ 0.72 2.06
+ 0.72 2.07
+ 0.72 2.08
+ 0.72 2.09
+ 0.72 2.1
+ 0.72 2.11
+ 0.72 2.12
+ 0.72 2.13
+ 0.72 2.14
+ 0.72 2.15
+ 0.72 2.16
+ 0.72 2.17
+ 0.72 2.18
+ 0.72 2.19
+ 0.72 2.2
+ 0.72 2.21
+ 0.72 2.22
+ 0.72 2.23
+ 0.72 2.24
+ 0.72 2.25
+ 0.72 2.26
+ 0.72 2.27
+ 0.72 2.28
+ 0.72 2.29
+ 0.72 2.3
+ 0.72 2.31
+ 0.72 2.32
+ 0.72 2.33
+ 0.72 2.34
+ 0.72 2.35
+ 0.72 2.36
+ 0.72 2.37
+ 0.72 2.38
+ 0.72 2.39
+ 0.72 2.4
+ 0.72 2.41
+ 0.72 2.42
+ 0.72 2.43
+ 0.72 2.44
+ 0.72 2.45
+ 0.72 2.46
+ 0.72 2.47
+ 0.72 2.48
+ 0.72 2.49
+ 0.72 2.5
+ 0.73 1.25
+ 0.73 1.26
+ 0.73 1.27
+ 0.73 1.28
+ 0.73 1.29
+ 0.73 1.3
+ 0.73 1.31
+ 0.73 1.32
+ 0.73 1.33
+ 0.73 1.34
+ 0.73 1.35
+ 0.73 1.36
+ 0.73 1.37
+ 0.73 1.38
+ 0.73 1.39
+ 0.73 1.4
+ 0.73 1.41
+ 0.73 1.42
+ 0.73 1.43
+ 0.73 1.44
+ 0.73 1.45
+ 0.73 1.46
+ 0.73 1.47
+ 0.73 1.48
+ 0.73 1.49
+ 0.73 1.5
+ 0.73 1.51
+ 0.73 1.52
+ 0.73 1.53
+ 0.73 1.54
+ 0.73 1.55
+ 0.73 1.56
+ 0.73 1.57
+ 0.73 1.58
+ 0.73 1.59
+ 0.73 1.6
+ 0.73 1.61
+ 0.73 1.62
+ 0.73 1.63
+ 0.73 1.64
+ 0.73 1.65
+ 0.73 1.66
+ 0.73 1.67
+ 0.73 1.68
+ 0.73 1.69
+ 0.73 1.7
+ 0.73 1.71
+ 0.73 1.72
+ 0.73 1.73
+ 0.73 1.74
+ 0.73 1.75
+ 0.73 1.76
+ 0.73 1.77
+ 0.73 1.78
+ 0.73 1.79
+ 0.73 1.8
+ 0.73 1.81
+ 0.73 1.82
+ 0.73 1.83
+ 0.73 1.84
+ 0.73 1.85
+ 0.73 1.86
+ 0.73 1.87
+ 0.73 1.88
+ 0.73 1.89
+ 0.73 1.9
+ 0.73 1.91
+ 0.73 1.92
+ 0.73 1.93
+ 0.73 1.94
+ 0.73 1.95
+ 0.73 1.96
+ 0.73 1.97
+ 0.73 1.98
+ 0.73 1.99
+ 0.73 2.0
+ 0.73 2.01
+ 0.73 2.02
+ 0.73 2.03
+ 0.73 2.04
+ 0.73 2.05
+ 0.73 2.06
+ 0.73 2.07
+ 0.73 2.08
+ 0.73 2.09
+ 0.73 2.1
+ 0.73 2.11
+ 0.73 2.12
+ 0.73 2.13
+ 0.73 2.14
+ 0.73 2.15
+ 0.73 2.16
+ 0.73 2.17
+ 0.73 2.18
+ 0.73 2.19
+ 0.73 2.2
+ 0.73 2.21
+ 0.73 2.22
+ 0.73 2.23
+ 0.73 2.24
+ 0.73 2.25
+ 0.73 2.26
+ 0.73 2.27
+ 0.73 2.28
+ 0.73 2.29
+ 0.73 2.3
+ 0.73 2.31
+ 0.73 2.32
+ 0.73 2.33
+ 0.73 2.34
+ 0.73 2.35
+ 0.73 2.36
+ 0.73 2.37
+ 0.73 2.38
+ 0.73 2.39
+ 0.73 2.4
+ 0.73 2.41
+ 0.73 2.42
+ 0.73 2.43
+ 0.73 2.44
+ 0.73 2.45
+ 0.73 2.46
+ 0.73 2.47
+ 0.73 2.48
+ 0.73 2.49
+ 0.73 2.5
+ 0.74 1.25
+ 0.74 1.26
+ 0.74 1.27
+ 0.74 1.28
+ 0.74 1.29
+ 0.74 1.3
+ 0.74 1.31
+ 0.74 1.32
+ 0.74 1.33
+ 0.74 1.34
+ 0.74 1.35
+ 0.74 1.36
+ 0.74 1.37
+ 0.74 1.38
+ 0.74 1.39
+ 0.74 1.4
+ 0.74 1.41
+ 0.74 1.42
+ 0.74 1.43
+ 0.74 1.44
+ 0.74 1.45
+ 0.74 1.46
+ 0.74 1.47
+ 0.74 1.48
+ 0.74 1.49
+ 0.74 1.5
+ 0.74 1.51
+ 0.74 1.52
+ 0.74 1.53
+ 0.74 1.54
+ 0.74 1.55
+ 0.74 1.56
+ 0.74 1.57
+ 0.74 1.58
+ 0.74 1.59
+ 0.74 1.6
+ 0.74 1.61
+ 0.74 1.62
+ 0.74 1.63
+ 0.74 1.64
+ 0.74 1.65
+ 0.74 1.66
+ 0.74 1.67
+ 0.74 1.68
+ 0.74 1.69
+ 0.74 1.7
+ 0.74 1.71
+ 0.74 1.72
+ 0.74 1.73
+ 0.74 1.74
+ 0.74 1.75
+ 0.74 1.76
+ 0.74 1.77
+ 0.74 1.78
+ 0.74 1.79
+ 0.74 1.8
+ 0.74 1.81
+ 0.74 1.82
+ 0.74 1.83
+ 0.74 1.84
+ 0.74 1.85
+ 0.74 1.86
+ 0.74 1.87
+ 0.74 1.88
+ 0.74 1.89
+ 0.74 1.9
+ 0.74 1.91
+ 0.74 1.92
+ 0.74 1.93
+ 0.74 1.94
+ 0.74 1.95
+ 0.74 1.96
+ 0.74 1.97
+ 0.74 1.98
+ 0.74 1.99
+ 0.74 2.0
+ 0.74 2.01
+ 0.74 2.02
+ 0.74 2.03
+ 0.74 2.04
+ 0.74 2.05
+ 0.74 2.06
+ 0.74 2.07
+ 0.74 2.08
+ 0.74 2.09
+ 0.74 2.1
+ 0.74 2.11
+ 0.74 2.12
+ 0.74 2.13
+ 0.74 2.14
+ 0.74 2.15
+ 0.74 2.16
+ 0.74 2.17
+ 0.74 2.18
+ 0.74 2.19
+ 0.74 2.2
+ 0.74 2.21
+ 0.74 2.22
+ 0.74 2.23
+ 0.74 2.24
+ 0.74 2.25
+ 0.74 2.26
+ 0.74 2.27
+ 0.74 2.28
+ 0.74 2.29
+ 0.74 2.3
+ 0.74 2.31
+ 0.74 2.32
+ 0.74 2.33
+ 0.74 2.34
+ 0.74 2.35
+ 0.74 2.36
+ 0.74 2.37
+ 0.74 2.38
+ 0.74 2.39
+ 0.74 2.4
+ 0.74 2.41
+ 0.74 2.42
+ 0.74 2.43
+ 0.74 2.44
+ 0.74 2.45
+ 0.74 2.46
+ 0.74 2.47
+ 0.74 2.48
+ 0.74 2.49
+ 0.74 2.5
+ 0.75 1.25
+ 0.75 1.26
+ 0.75 1.27
+ 0.75 1.28
+ 0.75 1.29
+ 0.75 1.3
+ 0.75 1.31
+ 0.75 1.32
+ 0.75 1.33
+ 0.75 1.34
+ 0.75 1.35
+ 0.75 1.36
+ 0.75 1.37
+ 0.75 1.38
+ 0.75 1.39
+ 0.75 1.4
+ 0.75 1.41
+ 0.75 1.42
+ 0.75 1.43
+ 0.75 1.44
+ 0.75 1.45
+ 0.75 1.46
+ 0.75 1.47
+ 0.75 1.48
+ 0.75 1.49
+ 0.75 1.5
+ 0.75 1.51
+ 0.75 1.52
+ 0.75 1.53
+ 0.75 1.54
+ 0.75 1.55
+ 0.75 1.56
+ 0.75 1.57
+ 0.75 1.58
+ 0.75 1.59
+ 0.75 1.6
+ 0.75 1.61
+ 0.75 1.62
+ 0.75 1.63
+ 0.75 1.64
+ 0.75 1.65
+ 0.75 1.66
+ 0.75 1.67
+ 0.75 1.68
+ 0.75 1.69
+ 0.75 1.7
+ 0.75 1.71
+ 0.75 1.72
+ 0.75 1.73
+ 0.75 1.74
+ 0.75 1.75
+ 0.75 1.76
+ 0.75 1.77
+ 0.75 1.78
+ 0.75 1.79
+ 0.75 1.8
+ 0.75 1.81
+ 0.75 1.82
+ 0.75 1.83
+ 0.75 1.84
+ 0.75 1.85
+ 0.75 1.86
+ 0.75 1.87
+ 0.75 1.88
+ 0.75 1.89
+ 0.75 1.9
+ 0.75 1.91
+ 0.75 1.92
+ 0.75 1.93
+ 0.75 1.94
+ 0.75 1.95
+ 0.75 1.96
+ 0.75 1.97
+ 0.75 1.98
+ 0.75 1.99
+ 0.75 2.0
+ 0.75 2.01
+ 0.75 2.02
+ 0.75 2.03
+ 0.75 2.04
+ 0.75 2.05
+ 0.75 2.06
+ 0.75 2.07
+ 0.75 2.08
+ 0.75 2.09
+ 0.75 2.1
+ 0.75 2.11
+ 0.75 2.12
+ 0.75 2.13
+ 0.75 2.14
+ 0.75 2.15
+ 0.75 2.16
+ 0.75 2.17
+ 0.75 2.18
+ 0.75 2.19
+ 0.75 2.2
+ 0.75 2.21
+ 0.75 2.22
+ 0.75 2.23
+ 0.75 2.24
+ 0.75 2.25
+ 0.75 2.26
+ 0.75 2.27
+ 0.75 2.28
+ 0.75 2.29
+ 0.75 2.3
+ 0.75 2.31
+ 0.75 2.32
+ 0.75 2.33
+ 0.75 2.34
+ 0.75 2.35
+ 0.75 2.36
+ 0.75 2.37
+ 0.75 2.38
+ 0.75 2.39
+ 0.75 2.4
+ 0.75 2.41
+ 0.75 2.42
+ 0.75 2.43
+ 0.75 2.44
+ 0.75 2.45
+ 0.75 2.46
+ 0.75 2.47
+ 0.75 2.48
+ 0.75 2.49
+ 0.75 2.5
+ 0.76 1.25
+ 0.76 1.26
+ 0.76 1.27
+ 0.76 1.28
+ 0.76 1.29
+ 0.76 1.3
+ 0.76 1.31
+ 0.76 1.32
+ 0.76 1.33
+ 0.76 1.34
+ 0.76 1.35
+ 0.76 1.36
+ 0.76 1.37
+ 0.76 1.38
+ 0.76 1.39
+ 0.76 1.4
+ 0.76 1.41
+ 0.76 1.42
+ 0.76 1.43
+ 0.76 1.44
+ 0.76 1.45
+ 0.76 1.46
+ 0.76 1.47
+ 0.76 1.48
+ 0.76 1.49
+ 0.76 1.5
+ 0.76 1.51
+ 0.76 1.52
+ 0.76 1.53
+ 0.76 1.54
+ 0.76 1.55
+ 0.76 1.56
+ 0.76 1.57
+ 0.76 1.58
+ 0.76 1.59
+ 0.76 1.6
+ 0.76 1.61
+ 0.76 1.62
+ 0.76 1.63
+ 0.76 1.64
+ 0.76 1.65
+ 0.76 1.66
+ 0.76 1.67
+ 0.76 1.68
+ 0.76 1.69
+ 0.76 1.7
+ 0.76 1.71
+ 0.76 1.72
+ 0.76 1.73
+ 0.76 1.74
+ 0.76 1.75
+ 0.76 1.76
+ 0.76 1.77
+ 0.76 1.78
+ 0.76 1.79
+ 0.76 1.8
+ 0.76 1.81
+ 0.76 1.82
+ 0.76 1.83
+ 0.76 1.84
+ 0.76 1.85
+ 0.76 1.86
+ 0.76 1.87
+ 0.76 1.88
+ 0.76 1.89
+ 0.76 1.9
+ 0.76 1.91
+ 0.76 1.92
+ 0.76 1.93
+ 0.76 1.94
+ 0.76 1.95
+ 0.76 1.96
+ 0.76 1.97
+ 0.76 1.98
+ 0.76 1.99
+ 0.76 2.0
+ 0.76 2.01
+ 0.76 2.02
+ 0.76 2.03
+ 0.76 2.04
+ 0.76 2.05
+ 0.76 2.06
+ 0.76 2.07
+ 0.76 2.08
+ 0.76 2.09
+ 0.76 2.1
+ 0.76 2.11
+ 0.76 2.12
+ 0.76 2.13
+ 0.76 2.14
+ 0.76 2.15
+ 0.76 2.16
+ 0.76 2.17
+ 0.76 2.18
+ 0.76 2.19
+ 0.76 2.2
+ 0.76 2.21
+ 0.76 2.22
+ 0.76 2.23
+ 0.76 2.24
+ 0.76 2.25
+ 0.76 2.26
+ 0.76 2.27
+ 0.76 2.28
+ 0.76 2.29
+ 0.76 2.3
+ 0.76 2.31
+ 0.76 2.32
+ 0.76 2.33
+ 0.76 2.34
+ 0.76 2.35
+ 0.76 2.36
+ 0.76 2.37
+ 0.76 2.38
+ 0.76 2.39
+ 0.76 2.4
+ 0.76 2.41
+ 0.76 2.42
+ 0.76 2.43
+ 0.76 2.44
+ 0.76 2.45
+ 0.76 2.46
+ 0.76 2.47
+ 0.76 2.48
+ 0.76 2.49
+ 0.76 2.5
+ 0.77 1.25
+ 0.77 1.26
+ 0.77 1.27
+ 0.77 1.28
+ 0.77 1.29
+ 0.77 1.3
+ 0.77 1.31
+ 0.77 1.32
+ 0.77 1.33
+ 0.77 1.34
+ 0.77 1.35
+ 0.77 1.36
+ 0.77 1.37
+ 0.77 1.38
+ 0.77 1.39
+ 0.77 1.4
+ 0.77 1.41
+ 0.77 1.42
+ 0.77 1.43
+ 0.77 1.44
+ 0.77 1.45
+ 0.77 1.46
+ 0.77 1.47
+ 0.77 1.48
+ 0.77 1.49
+ 0.77 1.5
+ 0.77 1.51
+ 0.77 1.52
+ 0.77 1.53
+ 0.77 1.54
+ 0.77 1.55
+ 0.77 1.56
+ 0.77 1.57
+ 0.77 1.58
+ 0.77 1.59
+ 0.77 1.6
+ 0.77 1.61
+ 0.77 1.62
+ 0.77 1.63
+ 0.77 1.64
+ 0.77 1.65
+ 0.77 1.66
+ 0.77 1.67
+ 0.77 1.68
+ 0.77 1.69
+ 0.77 1.7
+ 0.77 1.71
+ 0.77 1.72
+ 0.77 1.73
+ 0.77 1.74
+ 0.77 1.75
+ 0.77 1.76
+ 0.77 1.77
+ 0.77 1.78
+ 0.77 1.79
+ 0.77 1.8
+ 0.77 1.81
+ 0.77 1.82
+ 0.77 1.83
+ 0.77 1.84
+ 0.77 1.85
+ 0.77 1.86
+ 0.77 1.87
+ 0.77 1.88
+ 0.77 1.89
+ 0.77 1.9
+ 0.77 1.91
+ 0.77 1.92
+ 0.77 1.93
+ 0.77 1.94
+ 0.77 1.95
+ 0.77 1.96
+ 0.77 1.97
+ 0.77 1.98
+ 0.77 1.99
+ 0.77 2.0
+ 0.77 2.01
+ 0.77 2.02
+ 0.77 2.03
+ 0.77 2.04
+ 0.77 2.05
+ 0.77 2.06
+ 0.77 2.07
+ 0.77 2.08
+ 0.77 2.09
+ 0.77 2.1
+ 0.77 2.11
+ 0.77 2.12
+ 0.77 2.13
+ 0.77 2.14
+ 0.77 2.15
+ 0.77 2.16
+ 0.77 2.17
+ 0.77 2.18
+ 0.77 2.19
+ 0.77 2.2
+ 0.77 2.21
+ 0.77 2.22
+ 0.77 2.23
+ 0.77 2.24
+ 0.77 2.25
+ 0.77 2.26
+ 0.77 2.27
+ 0.77 2.28
+ 0.77 2.29
+ 0.77 2.3
+ 0.77 2.31
+ 0.77 2.32
+ 0.77 2.33
+ 0.77 2.34
+ 0.77 2.35
+ 0.77 2.36
+ 0.77 2.37
+ 0.77 2.38
+ 0.77 2.39
+ 0.77 2.4
+ 0.77 2.41
+ 0.77 2.42
+ 0.77 2.43
+ 0.77 2.44
+ 0.77 2.45
+ 0.77 2.46
+ 0.77 2.47
+ 0.77 2.48
+ 0.77 2.49
+ 0.77 2.5
+ 0.78 1.25
+ 0.78 1.26
+ 0.78 1.27
+ 0.78 1.28
+ 0.78 1.29
+ 0.78 1.3
+ 0.78 1.31
+ 0.78 1.32
+ 0.78 1.33
+ 0.78 1.34
+ 0.78 1.35
+ 0.78 1.36
+ 0.78 1.37
+ 0.78 1.38
+ 0.78 1.39
+ 0.78 1.4
+ 0.78 1.41
+ 0.78 1.42
+ 0.78 1.43
+ 0.78 1.44
+ 0.78 1.45
+ 0.78 1.46
+ 0.78 1.47
+ 0.78 1.48
+ 0.78 1.49
+ 0.78 1.5
+ 0.78 1.51
+ 0.78 1.52
+ 0.78 1.53
+ 0.78 1.54
+ 0.78 1.55
+ 0.78 1.56
+ 0.78 1.57
+ 0.78 1.58
+ 0.78 1.59
+ 0.78 1.6
+ 0.78 1.61
+ 0.78 1.62
+ 0.78 1.63
+ 0.78 1.64
+ 0.78 1.65
+ 0.78 1.66
+ 0.78 1.67
+ 0.78 1.68
+ 0.78 1.69
+ 0.78 1.7
+ 0.78 1.71
+ 0.78 1.72
+ 0.78 1.73
+ 0.78 1.74
+ 0.78 1.75
+ 0.78 1.76
+ 0.78 1.77
+ 0.78 1.78
+ 0.78 1.79
+ 0.78 1.8
+ 0.78 1.81
+ 0.78 1.82
+ 0.78 1.83
+ 0.78 1.84
+ 0.78 1.85
+ 0.78 1.86
+ 0.78 1.87
+ 0.78 1.88
+ 0.78 1.89
+ 0.78 1.9
+ 0.78 1.91
+ 0.78 1.92
+ 0.78 1.93
+ 0.78 1.94
+ 0.78 1.95
+ 0.78 1.96
+ 0.78 1.97
+ 0.78 1.98
+ 0.78 1.99
+ 0.78 2.0
+ 0.78 2.01
+ 0.78 2.02
+ 0.78 2.03
+ 0.78 2.04
+ 0.78 2.05
+ 0.78 2.06
+ 0.78 2.07
+ 0.78 2.08
+ 0.78 2.09
+ 0.78 2.1
+ 0.78 2.11
+ 0.78 2.12
+ 0.78 2.13
+ 0.78 2.14
+ 0.78 2.15
+ 0.78 2.16
+ 0.78 2.17
+ 0.78 2.18
+ 0.78 2.19
+ 0.78 2.2
+ 0.78 2.21
+ 0.78 2.22
+ 0.78 2.23
+ 0.78 2.24
+ 0.78 2.25
+ 0.78 2.26
+ 0.78 2.27
+ 0.78 2.28
+ 0.78 2.29
+ 0.78 2.3
+ 0.78 2.31
+ 0.78 2.32
+ 0.78 2.33
+ 0.78 2.34
+ 0.78 2.35
+ 0.78 2.36
+ 0.78 2.37
+ 0.78 2.38
+ 0.78 2.39
+ 0.78 2.4
+ 0.78 2.41
+ 0.78 2.42
+ 0.78 2.43
+ 0.78 2.44
+ 0.78 2.45
+ 0.78 2.46
+ 0.78 2.47
+ 0.78 2.48
+ 0.78 2.49
+ 0.78 2.5
+ 0.79 1.25
+ 0.79 1.26
+ 0.79 1.27
+ 0.79 1.28
+ 0.79 1.29
+ 0.79 1.3
+ 0.79 1.31
+ 0.79 1.32
+ 0.79 1.33
+ 0.79 1.34
+ 0.79 1.35
+ 0.79 1.36
+ 0.79 1.37
+ 0.79 1.38
+ 0.79 1.39
+ 0.79 1.4
+ 0.79 1.41
+ 0.79 1.42
+ 0.79 1.43
+ 0.79 1.44
+ 0.79 1.45
+ 0.79 1.46
+ 0.79 1.47
+ 0.79 1.48
+ 0.79 1.49
+ 0.79 1.5
+ 0.79 1.51
+ 0.79 1.52
+ 0.79 1.53
+ 0.79 1.54
+ 0.79 1.55
+ 0.79 1.56
+ 0.79 1.57
+ 0.79 1.58
+ 0.79 1.59
+ 0.79 1.6
+ 0.79 1.61
+ 0.79 1.62
+ 0.79 1.63
+ 0.79 1.64
+ 0.79 1.65
+ 0.79 1.66
+ 0.79 1.67
+ 0.79 1.68
+ 0.79 1.69
+ 0.79 1.7
+ 0.79 1.71
+ 0.79 1.72
+ 0.79 1.73
+ 0.79 1.74
+ 0.79 1.75
+ 0.79 1.76
+ 0.79 1.77
+ 0.79 1.78
+ 0.79 1.79
+ 0.79 1.8
+ 0.79 1.81
+ 0.79 1.82
+ 0.79 1.83
+ 0.79 1.84
+ 0.79 1.85
+ 0.79 1.86
+ 0.79 1.87
+ 0.79 1.88
+ 0.79 1.89
+ 0.79 1.9
+ 0.79 1.91
+ 0.79 1.92
+ 0.79 1.93
+ 0.79 1.94
+ 0.79 1.95
+ 0.79 1.96
+ 0.79 1.97
+ 0.79 1.98
+ 0.79 1.99
+ 0.79 2.0
+ 0.79 2.01
+ 0.79 2.02
+ 0.79 2.03
+ 0.79 2.04
+ 0.79 2.05
+ 0.79 2.06
+ 0.79 2.07
+ 0.79 2.08
+ 0.79 2.09
+ 0.79 2.1
+ 0.79 2.11
+ 0.79 2.12
+ 0.79 2.13
+ 0.79 2.14
+ 0.79 2.15
+ 0.79 2.16
+ 0.79 2.17
+ 0.79 2.18
+ 0.79 2.19
+ 0.79 2.2
+ 0.79 2.21
+ 0.79 2.22
+ 0.79 2.23
+ 0.79 2.24
+ 0.79 2.25
+ 0.79 2.26
+ 0.79 2.27
+ 0.79 2.28
+ 0.79 2.29
+ 0.79 2.3
+ 0.79 2.31
+ 0.79 2.32
+ 0.79 2.33
+ 0.79 2.34
+ 0.79 2.35
+ 0.79 2.36
+ 0.79 2.37
+ 0.79 2.38
+ 0.79 2.39
+ 0.79 2.4
+ 0.79 2.41
+ 0.79 2.42
+ 0.79 2.43
+ 0.79 2.44
+ 0.79 2.45
+ 0.79 2.46
+ 0.79 2.47
+ 0.79 2.48
+ 0.79 2.49
+ 0.79 2.5
+ 0.8 1.25
+ 0.8 1.26
+ 0.8 1.27
+ 0.8 1.28
+ 0.8 1.29
+ 0.8 1.3
+ 0.8 1.31
+ 0.8 1.32
+ 0.8 1.33
+ 0.8 1.34
+ 0.8 1.35
+ 0.8 1.36
+ 0.8 1.37
+ 0.8 1.38
+ 0.8 1.39
+ 0.8 1.4
+ 0.8 1.41
+ 0.8 1.42
+ 0.8 1.43
+ 0.8 1.44
+ 0.8 1.45
+ 0.8 1.46
+ 0.8 1.47
+ 0.8 1.48
+ 0.8 1.49
+ 0.8 1.5
+ 0.8 1.51
+ 0.8 1.52
+ 0.8 1.53
+ 0.8 1.54
+ 0.8 1.55
+ 0.8 1.56
+ 0.8 1.57
+ 0.8 1.58
+ 0.8 1.59
+ 0.8 1.6
+ 0.8 1.61
+ 0.8 1.62
+ 0.8 1.63
+ 0.8 1.64
+ 0.8 1.65
+ 0.8 1.66
+ 0.8 1.67
+ 0.8 1.68
+ 0.8 1.69
+ 0.8 1.7
+ 0.8 1.71
+ 0.8 1.72
+ 0.8 1.73
+ 0.8 1.74
+ 0.8 1.75
+ 0.8 1.76
+ 0.8 1.77
+ 0.8 1.78
+ 0.8 1.79
+ 0.8 1.8
+ 0.8 1.81
+ 0.8 1.82
+ 0.8 1.83
+ 0.8 1.84
+ 0.8 1.85
+ 0.8 1.86
+ 0.8 1.87
+ 0.8 1.88
+ 0.8 1.89
+ 0.8 1.9
+ 0.8 1.91
+ 0.8 1.92
+ 0.8 1.93
+ 0.8 1.94
+ 0.8 1.95
+ 0.8 1.96
+ 0.8 1.97
+ 0.8 1.98
+ 0.8 1.99
+ 0.8 2.0
+ 0.8 2.01
+ 0.8 2.02
+ 0.8 2.03
+ 0.8 2.04
+ 0.8 2.05
+ 0.8 2.06
+ 0.8 2.07
+ 0.8 2.08
+ 0.8 2.09
+ 0.8 2.1
+ 0.8 2.11
+ 0.8 2.12
+ 0.8 2.13
+ 0.8 2.14
+ 0.8 2.15
+ 0.8 2.16
+ 0.8 2.17
+ 0.8 2.18
+ 0.8 2.19
+ 0.8 2.2
+ 0.8 2.21
+ 0.8 2.22
+ 0.8 2.23
+ 0.8 2.24
+ 0.8 2.25
+ 0.8 2.26
+ 0.8 2.27
+ 0.8 2.28
+ 0.8 2.29
+ 0.8 2.3
+ 0.8 2.31
+ 0.8 2.32
+ 0.8 2.33
+ 0.8 2.34
+ 0.8 2.35
+ 0.8 2.36
+ 0.8 2.37
+ 0.8 2.38
+ 0.8 2.39
+ 0.8 2.4
+ 0.8 2.41
+ 0.8 2.42
+ 0.8 2.43
+ 0.8 2.44
+ 0.8 2.45
+ 0.8 2.46
+ 0.8 2.47
+ 0.8 2.48
+ 0.8 2.49
+ 0.8 2.5
.ENDDATA
