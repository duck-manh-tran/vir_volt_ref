
.option MEASFORM=3
.option RUNLVL=4
.option MEASDGT=6
.param vdd=0.8
.param k1 = 0.4
.param k2 = 0.3
.param k3 = 0.25
.param v_cap1='vdd*r_cap*k1'
.param v_cap2='vdd*r_cap*k2'
.param v_cap3='vdd*r_cap*k3'

.ic v(vdis)='vdd+0.01'

.meas tran t_dis1 TRIG v(vdis) val='v_cap1' FALL=1 TARG v(vdis) val='vdd*0.25' FALL=1
.meas tran t_dis2 TRIG v(vdis) val='v_cap2' FALL=1 TARG v(vdis) val='vdd*0.25' FALL=1
.meas tran t_dis3 TRIG v(vdis) val='v_cap3' FALL=1 TARG v(vdis) val='vdd*0.25' FALL=1

.tran 1n 8m sweep DATA=input

.DATA input
+ temp_val vdd r_cap
+ 0 0.4 1.25
+ 0 0.4 1.275
+ 0 0.4 1.3
+ 0 0.4 1.325
+ 0 0.4 1.35
+ 0 0.4 1.375
+ 0 0.4 1.4
+ 0 0.4 1.425
+ 0 0.4 1.45
+ 0 0.4 1.475
+ 0 0.4 1.5
+ 0 0.4 1.525
+ 0 0.4 1.55
+ 0 0.4 1.575
+ 0 0.4 1.6
+ 0 0.4 1.625
+ 0 0.4 1.65
+ 0 0.4 1.675
+ 0 0.4 1.7
+ 0 0.4 1.725
+ 0 0.4 1.75
+ 0 0.4 1.775
+ 0 0.4 1.8
+ 0 0.4 1.825
+ 0 0.4 1.85
+ 0 0.4 1.875
+ 0 0.4 1.9
+ 0 0.4 1.925
+ 0 0.4 1.95
+ 0 0.4 1.975
+ 0 0.4 2.0
+ 0 0.4 2.025
+ 0 0.4 2.05
+ 0 0.4 2.075
+ 0 0.4 2.1
+ 0 0.4 2.125
+ 0 0.4 2.15
+ 0 0.4 2.175
+ 0 0.4 2.2
+ 0 0.4 2.225
+ 0 0.4 2.25
+ 0 0.4 2.275
+ 0 0.4 2.3
+ 0 0.4 2.325
+ 0 0.4 2.35
+ 0 0.4 2.375
+ 0 0.4 2.4
+ 0 0.4 2.425
+ 0 0.4 2.45
+ 0 0.4 2.475
+ 0 0.4 2.5
+ 2 0.4 1.25
+ 2 0.4 1.275
+ 2 0.4 1.3
+ 2 0.4 1.325
+ 2 0.4 1.35
+ 2 0.4 1.375
+ 2 0.4 1.4
+ 2 0.4 1.425
+ 2 0.4 1.45
+ 2 0.4 1.475
+ 2 0.4 1.5
+ 2 0.4 1.525
+ 2 0.4 1.55
+ 2 0.4 1.575
+ 2 0.4 1.6
+ 2 0.4 1.625
+ 2 0.4 1.65
+ 2 0.4 1.675
+ 2 0.4 1.7
+ 2 0.4 1.725
+ 2 0.4 1.75
+ 2 0.4 1.775
+ 2 0.4 1.8
+ 2 0.4 1.825
+ 2 0.4 1.85
+ 2 0.4 1.875
+ 2 0.4 1.9
+ 2 0.4 1.925
+ 2 0.4 1.95
+ 2 0.4 1.975
+ 2 0.4 2.0
+ 2 0.4 2.025
+ 2 0.4 2.05
+ 2 0.4 2.075
+ 2 0.4 2.1
+ 2 0.4 2.125
+ 2 0.4 2.15
+ 2 0.4 2.175
+ 2 0.4 2.2
+ 2 0.4 2.225
+ 2 0.4 2.25
+ 2 0.4 2.275
+ 2 0.4 2.3
+ 2 0.4 2.325
+ 2 0.4 2.35
+ 2 0.4 2.375
+ 2 0.4 2.4
+ 2 0.4 2.425
+ 2 0.4 2.45
+ 2 0.4 2.475
+ 2 0.4 2.5
+ 4 0.4 1.25
+ 4 0.4 1.275
+ 4 0.4 1.3
+ 4 0.4 1.325
+ 4 0.4 1.35
+ 4 0.4 1.375
+ 4 0.4 1.4
+ 4 0.4 1.425
+ 4 0.4 1.45
+ 4 0.4 1.475
+ 4 0.4 1.5
+ 4 0.4 1.525
+ 4 0.4 1.55
+ 4 0.4 1.575
+ 4 0.4 1.6
+ 4 0.4 1.625
+ 4 0.4 1.65
+ 4 0.4 1.675
+ 4 0.4 1.7
+ 4 0.4 1.725
+ 4 0.4 1.75
+ 4 0.4 1.775
+ 4 0.4 1.8
+ 4 0.4 1.825
+ 4 0.4 1.85
+ 4 0.4 1.875
+ 4 0.4 1.9
+ 4 0.4 1.925
+ 4 0.4 1.95
+ 4 0.4 1.975
+ 4 0.4 2.0
+ 4 0.4 2.025
+ 4 0.4 2.05
+ 4 0.4 2.075
+ 4 0.4 2.1
+ 4 0.4 2.125
+ 4 0.4 2.15
+ 4 0.4 2.175
+ 4 0.4 2.2
+ 4 0.4 2.225
+ 4 0.4 2.25
+ 4 0.4 2.275
+ 4 0.4 2.3
+ 4 0.4 2.325
+ 4 0.4 2.35
+ 4 0.4 2.375
+ 4 0.4 2.4
+ 4 0.4 2.425
+ 4 0.4 2.45
+ 4 0.4 2.475
+ 4 0.4 2.5
+ 6 0.4 1.25
+ 6 0.4 1.275
+ 6 0.4 1.3
+ 6 0.4 1.325
+ 6 0.4 1.35
+ 6 0.4 1.375
+ 6 0.4 1.4
+ 6 0.4 1.425
+ 6 0.4 1.45
+ 6 0.4 1.475
+ 6 0.4 1.5
+ 6 0.4 1.525
+ 6 0.4 1.55
+ 6 0.4 1.575
+ 6 0.4 1.6
+ 6 0.4 1.625
+ 6 0.4 1.65
+ 6 0.4 1.675
+ 6 0.4 1.7
+ 6 0.4 1.725
+ 6 0.4 1.75
+ 6 0.4 1.775
+ 6 0.4 1.8
+ 6 0.4 1.825
+ 6 0.4 1.85
+ 6 0.4 1.875
+ 6 0.4 1.9
+ 6 0.4 1.925
+ 6 0.4 1.95
+ 6 0.4 1.975
+ 6 0.4 2.0
+ 6 0.4 2.025
+ 6 0.4 2.05
+ 6 0.4 2.075
+ 6 0.4 2.1
+ 6 0.4 2.125
+ 6 0.4 2.15
+ 6 0.4 2.175
+ 6 0.4 2.2
+ 6 0.4 2.225
+ 6 0.4 2.25
+ 6 0.4 2.275
+ 6 0.4 2.3
+ 6 0.4 2.325
+ 6 0.4 2.35
+ 6 0.4 2.375
+ 6 0.4 2.4
+ 6 0.4 2.425
+ 6 0.4 2.45
+ 6 0.4 2.475
+ 6 0.4 2.5
+ 8 0.4 1.25
+ 8 0.4 1.275
+ 8 0.4 1.3
+ 8 0.4 1.325
+ 8 0.4 1.35
+ 8 0.4 1.375
+ 8 0.4 1.4
+ 8 0.4 1.425
+ 8 0.4 1.45
+ 8 0.4 1.475
+ 8 0.4 1.5
+ 8 0.4 1.525
+ 8 0.4 1.55
+ 8 0.4 1.575
+ 8 0.4 1.6
+ 8 0.4 1.625
+ 8 0.4 1.65
+ 8 0.4 1.675
+ 8 0.4 1.7
+ 8 0.4 1.725
+ 8 0.4 1.75
+ 8 0.4 1.775
+ 8 0.4 1.8
+ 8 0.4 1.825
+ 8 0.4 1.85
+ 8 0.4 1.875
+ 8 0.4 1.9
+ 8 0.4 1.925
+ 8 0.4 1.95
+ 8 0.4 1.975
+ 8 0.4 2.0
+ 8 0.4 2.025
+ 8 0.4 2.05
+ 8 0.4 2.075
+ 8 0.4 2.1
+ 8 0.4 2.125
+ 8 0.4 2.15
+ 8 0.4 2.175
+ 8 0.4 2.2
+ 8 0.4 2.225
+ 8 0.4 2.25
+ 8 0.4 2.275
+ 8 0.4 2.3
+ 8 0.4 2.325
+ 8 0.4 2.35
+ 8 0.4 2.375
+ 8 0.4 2.4
+ 8 0.4 2.425
+ 8 0.4 2.45
+ 8 0.4 2.475
+ 8 0.4 2.5
+ 10 0.4 1.25
+ 10 0.4 1.275
+ 10 0.4 1.3
+ 10 0.4 1.325
+ 10 0.4 1.35
+ 10 0.4 1.375
+ 10 0.4 1.4
+ 10 0.4 1.425
+ 10 0.4 1.45
+ 10 0.4 1.475
+ 10 0.4 1.5
+ 10 0.4 1.525
+ 10 0.4 1.55
+ 10 0.4 1.575
+ 10 0.4 1.6
+ 10 0.4 1.625
+ 10 0.4 1.65
+ 10 0.4 1.675
+ 10 0.4 1.7
+ 10 0.4 1.725
+ 10 0.4 1.75
+ 10 0.4 1.775
+ 10 0.4 1.8
+ 10 0.4 1.825
+ 10 0.4 1.85
+ 10 0.4 1.875
+ 10 0.4 1.9
+ 10 0.4 1.925
+ 10 0.4 1.95
+ 10 0.4 1.975
+ 10 0.4 2.0
+ 10 0.4 2.025
+ 10 0.4 2.05
+ 10 0.4 2.075
+ 10 0.4 2.1
+ 10 0.4 2.125
+ 10 0.4 2.15
+ 10 0.4 2.175
+ 10 0.4 2.2
+ 10 0.4 2.225
+ 10 0.4 2.25
+ 10 0.4 2.275
+ 10 0.4 2.3
+ 10 0.4 2.325
+ 10 0.4 2.35
+ 10 0.4 2.375
+ 10 0.4 2.4
+ 10 0.4 2.425
+ 10 0.4 2.45
+ 10 0.4 2.475
+ 10 0.4 2.5
+ 12 0.4 1.25
+ 12 0.4 1.275
+ 12 0.4 1.3
+ 12 0.4 1.325
+ 12 0.4 1.35
+ 12 0.4 1.375
+ 12 0.4 1.4
+ 12 0.4 1.425
+ 12 0.4 1.45
+ 12 0.4 1.475
+ 12 0.4 1.5
+ 12 0.4 1.525
+ 12 0.4 1.55
+ 12 0.4 1.575
+ 12 0.4 1.6
+ 12 0.4 1.625
+ 12 0.4 1.65
+ 12 0.4 1.675
+ 12 0.4 1.7
+ 12 0.4 1.725
+ 12 0.4 1.75
+ 12 0.4 1.775
+ 12 0.4 1.8
+ 12 0.4 1.825
+ 12 0.4 1.85
+ 12 0.4 1.875
+ 12 0.4 1.9
+ 12 0.4 1.925
+ 12 0.4 1.95
+ 12 0.4 1.975
+ 12 0.4 2.0
+ 12 0.4 2.025
+ 12 0.4 2.05
+ 12 0.4 2.075
+ 12 0.4 2.1
+ 12 0.4 2.125
+ 12 0.4 2.15
+ 12 0.4 2.175
+ 12 0.4 2.2
+ 12 0.4 2.225
+ 12 0.4 2.25
+ 12 0.4 2.275
+ 12 0.4 2.3
+ 12 0.4 2.325
+ 12 0.4 2.35
+ 12 0.4 2.375
+ 12 0.4 2.4
+ 12 0.4 2.425
+ 12 0.4 2.45
+ 12 0.4 2.475
+ 12 0.4 2.5
+ 14 0.4 1.25
+ 14 0.4 1.275
+ 14 0.4 1.3
+ 14 0.4 1.325
+ 14 0.4 1.35
+ 14 0.4 1.375
+ 14 0.4 1.4
+ 14 0.4 1.425
+ 14 0.4 1.45
+ 14 0.4 1.475
+ 14 0.4 1.5
+ 14 0.4 1.525
+ 14 0.4 1.55
+ 14 0.4 1.575
+ 14 0.4 1.6
+ 14 0.4 1.625
+ 14 0.4 1.65
+ 14 0.4 1.675
+ 14 0.4 1.7
+ 14 0.4 1.725
+ 14 0.4 1.75
+ 14 0.4 1.775
+ 14 0.4 1.8
+ 14 0.4 1.825
+ 14 0.4 1.85
+ 14 0.4 1.875
+ 14 0.4 1.9
+ 14 0.4 1.925
+ 14 0.4 1.95
+ 14 0.4 1.975
+ 14 0.4 2.0
+ 14 0.4 2.025
+ 14 0.4 2.05
+ 14 0.4 2.075
+ 14 0.4 2.1
+ 14 0.4 2.125
+ 14 0.4 2.15
+ 14 0.4 2.175
+ 14 0.4 2.2
+ 14 0.4 2.225
+ 14 0.4 2.25
+ 14 0.4 2.275
+ 14 0.4 2.3
+ 14 0.4 2.325
+ 14 0.4 2.35
+ 14 0.4 2.375
+ 14 0.4 2.4
+ 14 0.4 2.425
+ 14 0.4 2.45
+ 14 0.4 2.475
+ 14 0.4 2.5
+ 16 0.4 1.25
+ 16 0.4 1.275
+ 16 0.4 1.3
+ 16 0.4 1.325
+ 16 0.4 1.35
+ 16 0.4 1.375
+ 16 0.4 1.4
+ 16 0.4 1.425
+ 16 0.4 1.45
+ 16 0.4 1.475
+ 16 0.4 1.5
+ 16 0.4 1.525
+ 16 0.4 1.55
+ 16 0.4 1.575
+ 16 0.4 1.6
+ 16 0.4 1.625
+ 16 0.4 1.65
+ 16 0.4 1.675
+ 16 0.4 1.7
+ 16 0.4 1.725
+ 16 0.4 1.75
+ 16 0.4 1.775
+ 16 0.4 1.8
+ 16 0.4 1.825
+ 16 0.4 1.85
+ 16 0.4 1.875
+ 16 0.4 1.9
+ 16 0.4 1.925
+ 16 0.4 1.95
+ 16 0.4 1.975
+ 16 0.4 2.0
+ 16 0.4 2.025
+ 16 0.4 2.05
+ 16 0.4 2.075
+ 16 0.4 2.1
+ 16 0.4 2.125
+ 16 0.4 2.15
+ 16 0.4 2.175
+ 16 0.4 2.2
+ 16 0.4 2.225
+ 16 0.4 2.25
+ 16 0.4 2.275
+ 16 0.4 2.3
+ 16 0.4 2.325
+ 16 0.4 2.35
+ 16 0.4 2.375
+ 16 0.4 2.4
+ 16 0.4 2.425
+ 16 0.4 2.45
+ 16 0.4 2.475
+ 16 0.4 2.5
+ 18 0.4 1.25
+ 18 0.4 1.275
+ 18 0.4 1.3
+ 18 0.4 1.325
+ 18 0.4 1.35
+ 18 0.4 1.375
+ 18 0.4 1.4
+ 18 0.4 1.425
+ 18 0.4 1.45
+ 18 0.4 1.475
+ 18 0.4 1.5
+ 18 0.4 1.525
+ 18 0.4 1.55
+ 18 0.4 1.575
+ 18 0.4 1.6
+ 18 0.4 1.625
+ 18 0.4 1.65
+ 18 0.4 1.675
+ 18 0.4 1.7
+ 18 0.4 1.725
+ 18 0.4 1.75
+ 18 0.4 1.775
+ 18 0.4 1.8
+ 18 0.4 1.825
+ 18 0.4 1.85
+ 18 0.4 1.875
+ 18 0.4 1.9
+ 18 0.4 1.925
+ 18 0.4 1.95
+ 18 0.4 1.975
+ 18 0.4 2.0
+ 18 0.4 2.025
+ 18 0.4 2.05
+ 18 0.4 2.075
+ 18 0.4 2.1
+ 18 0.4 2.125
+ 18 0.4 2.15
+ 18 0.4 2.175
+ 18 0.4 2.2
+ 18 0.4 2.225
+ 18 0.4 2.25
+ 18 0.4 2.275
+ 18 0.4 2.3
+ 18 0.4 2.325
+ 18 0.4 2.35
+ 18 0.4 2.375
+ 18 0.4 2.4
+ 18 0.4 2.425
+ 18 0.4 2.45
+ 18 0.4 2.475
+ 18 0.4 2.5
+ 20 0.4 1.25
+ 20 0.4 1.275
+ 20 0.4 1.3
+ 20 0.4 1.325
+ 20 0.4 1.35
+ 20 0.4 1.375
+ 20 0.4 1.4
+ 20 0.4 1.425
+ 20 0.4 1.45
+ 20 0.4 1.475
+ 20 0.4 1.5
+ 20 0.4 1.525
+ 20 0.4 1.55
+ 20 0.4 1.575
+ 20 0.4 1.6
+ 20 0.4 1.625
+ 20 0.4 1.65
+ 20 0.4 1.675
+ 20 0.4 1.7
+ 20 0.4 1.725
+ 20 0.4 1.75
+ 20 0.4 1.775
+ 20 0.4 1.8
+ 20 0.4 1.825
+ 20 0.4 1.85
+ 20 0.4 1.875
+ 20 0.4 1.9
+ 20 0.4 1.925
+ 20 0.4 1.95
+ 20 0.4 1.975
+ 20 0.4 2.0
+ 20 0.4 2.025
+ 20 0.4 2.05
+ 20 0.4 2.075
+ 20 0.4 2.1
+ 20 0.4 2.125
+ 20 0.4 2.15
+ 20 0.4 2.175
+ 20 0.4 2.2
+ 20 0.4 2.225
+ 20 0.4 2.25
+ 20 0.4 2.275
+ 20 0.4 2.3
+ 20 0.4 2.325
+ 20 0.4 2.35
+ 20 0.4 2.375
+ 20 0.4 2.4
+ 20 0.4 2.425
+ 20 0.4 2.45
+ 20 0.4 2.475
+ 20 0.4 2.5
+ 22 0.4 1.25
+ 22 0.4 1.275
+ 22 0.4 1.3
+ 22 0.4 1.325
+ 22 0.4 1.35
+ 22 0.4 1.375
+ 22 0.4 1.4
+ 22 0.4 1.425
+ 22 0.4 1.45
+ 22 0.4 1.475
+ 22 0.4 1.5
+ 22 0.4 1.525
+ 22 0.4 1.55
+ 22 0.4 1.575
+ 22 0.4 1.6
+ 22 0.4 1.625
+ 22 0.4 1.65
+ 22 0.4 1.675
+ 22 0.4 1.7
+ 22 0.4 1.725
+ 22 0.4 1.75
+ 22 0.4 1.775
+ 22 0.4 1.8
+ 22 0.4 1.825
+ 22 0.4 1.85
+ 22 0.4 1.875
+ 22 0.4 1.9
+ 22 0.4 1.925
+ 22 0.4 1.95
+ 22 0.4 1.975
+ 22 0.4 2.0
+ 22 0.4 2.025
+ 22 0.4 2.05
+ 22 0.4 2.075
+ 22 0.4 2.1
+ 22 0.4 2.125
+ 22 0.4 2.15
+ 22 0.4 2.175
+ 22 0.4 2.2
+ 22 0.4 2.225
+ 22 0.4 2.25
+ 22 0.4 2.275
+ 22 0.4 2.3
+ 22 0.4 2.325
+ 22 0.4 2.35
+ 22 0.4 2.375
+ 22 0.4 2.4
+ 22 0.4 2.425
+ 22 0.4 2.45
+ 22 0.4 2.475
+ 22 0.4 2.5
+ 24 0.4 1.25
+ 24 0.4 1.275
+ 24 0.4 1.3
+ 24 0.4 1.325
+ 24 0.4 1.35
+ 24 0.4 1.375
+ 24 0.4 1.4
+ 24 0.4 1.425
+ 24 0.4 1.45
+ 24 0.4 1.475
+ 24 0.4 1.5
+ 24 0.4 1.525
+ 24 0.4 1.55
+ 24 0.4 1.575
+ 24 0.4 1.6
+ 24 0.4 1.625
+ 24 0.4 1.65
+ 24 0.4 1.675
+ 24 0.4 1.7
+ 24 0.4 1.725
+ 24 0.4 1.75
+ 24 0.4 1.775
+ 24 0.4 1.8
+ 24 0.4 1.825
+ 24 0.4 1.85
+ 24 0.4 1.875
+ 24 0.4 1.9
+ 24 0.4 1.925
+ 24 0.4 1.95
+ 24 0.4 1.975
+ 24 0.4 2.0
+ 24 0.4 2.025
+ 24 0.4 2.05
+ 24 0.4 2.075
+ 24 0.4 2.1
+ 24 0.4 2.125
+ 24 0.4 2.15
+ 24 0.4 2.175
+ 24 0.4 2.2
+ 24 0.4 2.225
+ 24 0.4 2.25
+ 24 0.4 2.275
+ 24 0.4 2.3
+ 24 0.4 2.325
+ 24 0.4 2.35
+ 24 0.4 2.375
+ 24 0.4 2.4
+ 24 0.4 2.425
+ 24 0.4 2.45
+ 24 0.4 2.475
+ 24 0.4 2.5
+ 26 0.4 1.25
+ 26 0.4 1.275
+ 26 0.4 1.3
+ 26 0.4 1.325
+ 26 0.4 1.35
+ 26 0.4 1.375
+ 26 0.4 1.4
+ 26 0.4 1.425
+ 26 0.4 1.45
+ 26 0.4 1.475
+ 26 0.4 1.5
+ 26 0.4 1.525
+ 26 0.4 1.55
+ 26 0.4 1.575
+ 26 0.4 1.6
+ 26 0.4 1.625
+ 26 0.4 1.65
+ 26 0.4 1.675
+ 26 0.4 1.7
+ 26 0.4 1.725
+ 26 0.4 1.75
+ 26 0.4 1.775
+ 26 0.4 1.8
+ 26 0.4 1.825
+ 26 0.4 1.85
+ 26 0.4 1.875
+ 26 0.4 1.9
+ 26 0.4 1.925
+ 26 0.4 1.95
+ 26 0.4 1.975
+ 26 0.4 2.0
+ 26 0.4 2.025
+ 26 0.4 2.05
+ 26 0.4 2.075
+ 26 0.4 2.1
+ 26 0.4 2.125
+ 26 0.4 2.15
+ 26 0.4 2.175
+ 26 0.4 2.2
+ 26 0.4 2.225
+ 26 0.4 2.25
+ 26 0.4 2.275
+ 26 0.4 2.3
+ 26 0.4 2.325
+ 26 0.4 2.35
+ 26 0.4 2.375
+ 26 0.4 2.4
+ 26 0.4 2.425
+ 26 0.4 2.45
+ 26 0.4 2.475
+ 26 0.4 2.5
+ 28 0.4 1.25
+ 28 0.4 1.275
+ 28 0.4 1.3
+ 28 0.4 1.325
+ 28 0.4 1.35
+ 28 0.4 1.375
+ 28 0.4 1.4
+ 28 0.4 1.425
+ 28 0.4 1.45
+ 28 0.4 1.475
+ 28 0.4 1.5
+ 28 0.4 1.525
+ 28 0.4 1.55
+ 28 0.4 1.575
+ 28 0.4 1.6
+ 28 0.4 1.625
+ 28 0.4 1.65
+ 28 0.4 1.675
+ 28 0.4 1.7
+ 28 0.4 1.725
+ 28 0.4 1.75
+ 28 0.4 1.775
+ 28 0.4 1.8
+ 28 0.4 1.825
+ 28 0.4 1.85
+ 28 0.4 1.875
+ 28 0.4 1.9
+ 28 0.4 1.925
+ 28 0.4 1.95
+ 28 0.4 1.975
+ 28 0.4 2.0
+ 28 0.4 2.025
+ 28 0.4 2.05
+ 28 0.4 2.075
+ 28 0.4 2.1
+ 28 0.4 2.125
+ 28 0.4 2.15
+ 28 0.4 2.175
+ 28 0.4 2.2
+ 28 0.4 2.225
+ 28 0.4 2.25
+ 28 0.4 2.275
+ 28 0.4 2.3
+ 28 0.4 2.325
+ 28 0.4 2.35
+ 28 0.4 2.375
+ 28 0.4 2.4
+ 28 0.4 2.425
+ 28 0.4 2.45
+ 28 0.4 2.475
+ 28 0.4 2.5
+ 30 0.4 1.25
+ 30 0.4 1.275
+ 30 0.4 1.3
+ 30 0.4 1.325
+ 30 0.4 1.35
+ 30 0.4 1.375
+ 30 0.4 1.4
+ 30 0.4 1.425
+ 30 0.4 1.45
+ 30 0.4 1.475
+ 30 0.4 1.5
+ 30 0.4 1.525
+ 30 0.4 1.55
+ 30 0.4 1.575
+ 30 0.4 1.6
+ 30 0.4 1.625
+ 30 0.4 1.65
+ 30 0.4 1.675
+ 30 0.4 1.7
+ 30 0.4 1.725
+ 30 0.4 1.75
+ 30 0.4 1.775
+ 30 0.4 1.8
+ 30 0.4 1.825
+ 30 0.4 1.85
+ 30 0.4 1.875
+ 30 0.4 1.9
+ 30 0.4 1.925
+ 30 0.4 1.95
+ 30 0.4 1.975
+ 30 0.4 2.0
+ 30 0.4 2.025
+ 30 0.4 2.05
+ 30 0.4 2.075
+ 30 0.4 2.1
+ 30 0.4 2.125
+ 30 0.4 2.15
+ 30 0.4 2.175
+ 30 0.4 2.2
+ 30 0.4 2.225
+ 30 0.4 2.25
+ 30 0.4 2.275
+ 30 0.4 2.3
+ 30 0.4 2.325
+ 30 0.4 2.35
+ 30 0.4 2.375
+ 30 0.4 2.4
+ 30 0.4 2.425
+ 30 0.4 2.45
+ 30 0.4 2.475
+ 30 0.4 2.5
+ 32 0.4 1.25
+ 32 0.4 1.275
+ 32 0.4 1.3
+ 32 0.4 1.325
+ 32 0.4 1.35
+ 32 0.4 1.375
+ 32 0.4 1.4
+ 32 0.4 1.425
+ 32 0.4 1.45
+ 32 0.4 1.475
+ 32 0.4 1.5
+ 32 0.4 1.525
+ 32 0.4 1.55
+ 32 0.4 1.575
+ 32 0.4 1.6
+ 32 0.4 1.625
+ 32 0.4 1.65
+ 32 0.4 1.675
+ 32 0.4 1.7
+ 32 0.4 1.725
+ 32 0.4 1.75
+ 32 0.4 1.775
+ 32 0.4 1.8
+ 32 0.4 1.825
+ 32 0.4 1.85
+ 32 0.4 1.875
+ 32 0.4 1.9
+ 32 0.4 1.925
+ 32 0.4 1.95
+ 32 0.4 1.975
+ 32 0.4 2.0
+ 32 0.4 2.025
+ 32 0.4 2.05
+ 32 0.4 2.075
+ 32 0.4 2.1
+ 32 0.4 2.125
+ 32 0.4 2.15
+ 32 0.4 2.175
+ 32 0.4 2.2
+ 32 0.4 2.225
+ 32 0.4 2.25
+ 32 0.4 2.275
+ 32 0.4 2.3
+ 32 0.4 2.325
+ 32 0.4 2.35
+ 32 0.4 2.375
+ 32 0.4 2.4
+ 32 0.4 2.425
+ 32 0.4 2.45
+ 32 0.4 2.475
+ 32 0.4 2.5
+ 34 0.4 1.25
+ 34 0.4 1.275
+ 34 0.4 1.3
+ 34 0.4 1.325
+ 34 0.4 1.35
+ 34 0.4 1.375
+ 34 0.4 1.4
+ 34 0.4 1.425
+ 34 0.4 1.45
+ 34 0.4 1.475
+ 34 0.4 1.5
+ 34 0.4 1.525
+ 34 0.4 1.55
+ 34 0.4 1.575
+ 34 0.4 1.6
+ 34 0.4 1.625
+ 34 0.4 1.65
+ 34 0.4 1.675
+ 34 0.4 1.7
+ 34 0.4 1.725
+ 34 0.4 1.75
+ 34 0.4 1.775
+ 34 0.4 1.8
+ 34 0.4 1.825
+ 34 0.4 1.85
+ 34 0.4 1.875
+ 34 0.4 1.9
+ 34 0.4 1.925
+ 34 0.4 1.95
+ 34 0.4 1.975
+ 34 0.4 2.0
+ 34 0.4 2.025
+ 34 0.4 2.05
+ 34 0.4 2.075
+ 34 0.4 2.1
+ 34 0.4 2.125
+ 34 0.4 2.15
+ 34 0.4 2.175
+ 34 0.4 2.2
+ 34 0.4 2.225
+ 34 0.4 2.25
+ 34 0.4 2.275
+ 34 0.4 2.3
+ 34 0.4 2.325
+ 34 0.4 2.35
+ 34 0.4 2.375
+ 34 0.4 2.4
+ 34 0.4 2.425
+ 34 0.4 2.45
+ 34 0.4 2.475
+ 34 0.4 2.5
+ 36 0.4 1.25
+ 36 0.4 1.275
+ 36 0.4 1.3
+ 36 0.4 1.325
+ 36 0.4 1.35
+ 36 0.4 1.375
+ 36 0.4 1.4
+ 36 0.4 1.425
+ 36 0.4 1.45
+ 36 0.4 1.475
+ 36 0.4 1.5
+ 36 0.4 1.525
+ 36 0.4 1.55
+ 36 0.4 1.575
+ 36 0.4 1.6
+ 36 0.4 1.625
+ 36 0.4 1.65
+ 36 0.4 1.675
+ 36 0.4 1.7
+ 36 0.4 1.725
+ 36 0.4 1.75
+ 36 0.4 1.775
+ 36 0.4 1.8
+ 36 0.4 1.825
+ 36 0.4 1.85
+ 36 0.4 1.875
+ 36 0.4 1.9
+ 36 0.4 1.925
+ 36 0.4 1.95
+ 36 0.4 1.975
+ 36 0.4 2.0
+ 36 0.4 2.025
+ 36 0.4 2.05
+ 36 0.4 2.075
+ 36 0.4 2.1
+ 36 0.4 2.125
+ 36 0.4 2.15
+ 36 0.4 2.175
+ 36 0.4 2.2
+ 36 0.4 2.225
+ 36 0.4 2.25
+ 36 0.4 2.275
+ 36 0.4 2.3
+ 36 0.4 2.325
+ 36 0.4 2.35
+ 36 0.4 2.375
+ 36 0.4 2.4
+ 36 0.4 2.425
+ 36 0.4 2.45
+ 36 0.4 2.475
+ 36 0.4 2.5
+ 38 0.4 1.25
+ 38 0.4 1.275
+ 38 0.4 1.3
+ 38 0.4 1.325
+ 38 0.4 1.35
+ 38 0.4 1.375
+ 38 0.4 1.4
+ 38 0.4 1.425
+ 38 0.4 1.45
+ 38 0.4 1.475
+ 38 0.4 1.5
+ 38 0.4 1.525
+ 38 0.4 1.55
+ 38 0.4 1.575
+ 38 0.4 1.6
+ 38 0.4 1.625
+ 38 0.4 1.65
+ 38 0.4 1.675
+ 38 0.4 1.7
+ 38 0.4 1.725
+ 38 0.4 1.75
+ 38 0.4 1.775
+ 38 0.4 1.8
+ 38 0.4 1.825
+ 38 0.4 1.85
+ 38 0.4 1.875
+ 38 0.4 1.9
+ 38 0.4 1.925
+ 38 0.4 1.95
+ 38 0.4 1.975
+ 38 0.4 2.0
+ 38 0.4 2.025
+ 38 0.4 2.05
+ 38 0.4 2.075
+ 38 0.4 2.1
+ 38 0.4 2.125
+ 38 0.4 2.15
+ 38 0.4 2.175
+ 38 0.4 2.2
+ 38 0.4 2.225
+ 38 0.4 2.25
+ 38 0.4 2.275
+ 38 0.4 2.3
+ 38 0.4 2.325
+ 38 0.4 2.35
+ 38 0.4 2.375
+ 38 0.4 2.4
+ 38 0.4 2.425
+ 38 0.4 2.45
+ 38 0.4 2.475
+ 38 0.4 2.5
+ 40 0.4 1.25
+ 40 0.4 1.275
+ 40 0.4 1.3
+ 40 0.4 1.325
+ 40 0.4 1.35
+ 40 0.4 1.375
+ 40 0.4 1.4
+ 40 0.4 1.425
+ 40 0.4 1.45
+ 40 0.4 1.475
+ 40 0.4 1.5
+ 40 0.4 1.525
+ 40 0.4 1.55
+ 40 0.4 1.575
+ 40 0.4 1.6
+ 40 0.4 1.625
+ 40 0.4 1.65
+ 40 0.4 1.675
+ 40 0.4 1.7
+ 40 0.4 1.725
+ 40 0.4 1.75
+ 40 0.4 1.775
+ 40 0.4 1.8
+ 40 0.4 1.825
+ 40 0.4 1.85
+ 40 0.4 1.875
+ 40 0.4 1.9
+ 40 0.4 1.925
+ 40 0.4 1.95
+ 40 0.4 1.975
+ 40 0.4 2.0
+ 40 0.4 2.025
+ 40 0.4 2.05
+ 40 0.4 2.075
+ 40 0.4 2.1
+ 40 0.4 2.125
+ 40 0.4 2.15
+ 40 0.4 2.175
+ 40 0.4 2.2
+ 40 0.4 2.225
+ 40 0.4 2.25
+ 40 0.4 2.275
+ 40 0.4 2.3
+ 40 0.4 2.325
+ 40 0.4 2.35
+ 40 0.4 2.375
+ 40 0.4 2.4
+ 40 0.4 2.425
+ 40 0.4 2.45
+ 40 0.4 2.475
+ 40 0.4 2.5
+ 42 0.4 1.25
+ 42 0.4 1.275
+ 42 0.4 1.3
+ 42 0.4 1.325
+ 42 0.4 1.35
+ 42 0.4 1.375
+ 42 0.4 1.4
+ 42 0.4 1.425
+ 42 0.4 1.45
+ 42 0.4 1.475
+ 42 0.4 1.5
+ 42 0.4 1.525
+ 42 0.4 1.55
+ 42 0.4 1.575
+ 42 0.4 1.6
+ 42 0.4 1.625
+ 42 0.4 1.65
+ 42 0.4 1.675
+ 42 0.4 1.7
+ 42 0.4 1.725
+ 42 0.4 1.75
+ 42 0.4 1.775
+ 42 0.4 1.8
+ 42 0.4 1.825
+ 42 0.4 1.85
+ 42 0.4 1.875
+ 42 0.4 1.9
+ 42 0.4 1.925
+ 42 0.4 1.95
+ 42 0.4 1.975
+ 42 0.4 2.0
+ 42 0.4 2.025
+ 42 0.4 2.05
+ 42 0.4 2.075
+ 42 0.4 2.1
+ 42 0.4 2.125
+ 42 0.4 2.15
+ 42 0.4 2.175
+ 42 0.4 2.2
+ 42 0.4 2.225
+ 42 0.4 2.25
+ 42 0.4 2.275
+ 42 0.4 2.3
+ 42 0.4 2.325
+ 42 0.4 2.35
+ 42 0.4 2.375
+ 42 0.4 2.4
+ 42 0.4 2.425
+ 42 0.4 2.45
+ 42 0.4 2.475
+ 42 0.4 2.5
+ 44 0.4 1.25
+ 44 0.4 1.275
+ 44 0.4 1.3
+ 44 0.4 1.325
+ 44 0.4 1.35
+ 44 0.4 1.375
+ 44 0.4 1.4
+ 44 0.4 1.425
+ 44 0.4 1.45
+ 44 0.4 1.475
+ 44 0.4 1.5
+ 44 0.4 1.525
+ 44 0.4 1.55
+ 44 0.4 1.575
+ 44 0.4 1.6
+ 44 0.4 1.625
+ 44 0.4 1.65
+ 44 0.4 1.675
+ 44 0.4 1.7
+ 44 0.4 1.725
+ 44 0.4 1.75
+ 44 0.4 1.775
+ 44 0.4 1.8
+ 44 0.4 1.825
+ 44 0.4 1.85
+ 44 0.4 1.875
+ 44 0.4 1.9
+ 44 0.4 1.925
+ 44 0.4 1.95
+ 44 0.4 1.975
+ 44 0.4 2.0
+ 44 0.4 2.025
+ 44 0.4 2.05
+ 44 0.4 2.075
+ 44 0.4 2.1
+ 44 0.4 2.125
+ 44 0.4 2.15
+ 44 0.4 2.175
+ 44 0.4 2.2
+ 44 0.4 2.225
+ 44 0.4 2.25
+ 44 0.4 2.275
+ 44 0.4 2.3
+ 44 0.4 2.325
+ 44 0.4 2.35
+ 44 0.4 2.375
+ 44 0.4 2.4
+ 44 0.4 2.425
+ 44 0.4 2.45
+ 44 0.4 2.475
+ 44 0.4 2.5
+ 46 0.4 1.25
+ 46 0.4 1.275
+ 46 0.4 1.3
+ 46 0.4 1.325
+ 46 0.4 1.35
+ 46 0.4 1.375
+ 46 0.4 1.4
+ 46 0.4 1.425
+ 46 0.4 1.45
+ 46 0.4 1.475
+ 46 0.4 1.5
+ 46 0.4 1.525
+ 46 0.4 1.55
+ 46 0.4 1.575
+ 46 0.4 1.6
+ 46 0.4 1.625
+ 46 0.4 1.65
+ 46 0.4 1.675
+ 46 0.4 1.7
+ 46 0.4 1.725
+ 46 0.4 1.75
+ 46 0.4 1.775
+ 46 0.4 1.8
+ 46 0.4 1.825
+ 46 0.4 1.85
+ 46 0.4 1.875
+ 46 0.4 1.9
+ 46 0.4 1.925
+ 46 0.4 1.95
+ 46 0.4 1.975
+ 46 0.4 2.0
+ 46 0.4 2.025
+ 46 0.4 2.05
+ 46 0.4 2.075
+ 46 0.4 2.1
+ 46 0.4 2.125
+ 46 0.4 2.15
+ 46 0.4 2.175
+ 46 0.4 2.2
+ 46 0.4 2.225
+ 46 0.4 2.25
+ 46 0.4 2.275
+ 46 0.4 2.3
+ 46 0.4 2.325
+ 46 0.4 2.35
+ 46 0.4 2.375
+ 46 0.4 2.4
+ 46 0.4 2.425
+ 46 0.4 2.45
+ 46 0.4 2.475
+ 46 0.4 2.5
+ 48 0.4 1.25
+ 48 0.4 1.275
+ 48 0.4 1.3
+ 48 0.4 1.325
+ 48 0.4 1.35
+ 48 0.4 1.375
+ 48 0.4 1.4
+ 48 0.4 1.425
+ 48 0.4 1.45
+ 48 0.4 1.475
+ 48 0.4 1.5
+ 48 0.4 1.525
+ 48 0.4 1.55
+ 48 0.4 1.575
+ 48 0.4 1.6
+ 48 0.4 1.625
+ 48 0.4 1.65
+ 48 0.4 1.675
+ 48 0.4 1.7
+ 48 0.4 1.725
+ 48 0.4 1.75
+ 48 0.4 1.775
+ 48 0.4 1.8
+ 48 0.4 1.825
+ 48 0.4 1.85
+ 48 0.4 1.875
+ 48 0.4 1.9
+ 48 0.4 1.925
+ 48 0.4 1.95
+ 48 0.4 1.975
+ 48 0.4 2.0
+ 48 0.4 2.025
+ 48 0.4 2.05
+ 48 0.4 2.075
+ 48 0.4 2.1
+ 48 0.4 2.125
+ 48 0.4 2.15
+ 48 0.4 2.175
+ 48 0.4 2.2
+ 48 0.4 2.225
+ 48 0.4 2.25
+ 48 0.4 2.275
+ 48 0.4 2.3
+ 48 0.4 2.325
+ 48 0.4 2.35
+ 48 0.4 2.375
+ 48 0.4 2.4
+ 48 0.4 2.425
+ 48 0.4 2.45
+ 48 0.4 2.475
+ 48 0.4 2.5
+ 50 0.4 1.25
+ 50 0.4 1.275
+ 50 0.4 1.3
+ 50 0.4 1.325
+ 50 0.4 1.35
+ 50 0.4 1.375
+ 50 0.4 1.4
+ 50 0.4 1.425
+ 50 0.4 1.45
+ 50 0.4 1.475
+ 50 0.4 1.5
+ 50 0.4 1.525
+ 50 0.4 1.55
+ 50 0.4 1.575
+ 50 0.4 1.6
+ 50 0.4 1.625
+ 50 0.4 1.65
+ 50 0.4 1.675
+ 50 0.4 1.7
+ 50 0.4 1.725
+ 50 0.4 1.75
+ 50 0.4 1.775
+ 50 0.4 1.8
+ 50 0.4 1.825
+ 50 0.4 1.85
+ 50 0.4 1.875
+ 50 0.4 1.9
+ 50 0.4 1.925
+ 50 0.4 1.95
+ 50 0.4 1.975
+ 50 0.4 2.0
+ 50 0.4 2.025
+ 50 0.4 2.05
+ 50 0.4 2.075
+ 50 0.4 2.1
+ 50 0.4 2.125
+ 50 0.4 2.15
+ 50 0.4 2.175
+ 50 0.4 2.2
+ 50 0.4 2.225
+ 50 0.4 2.25
+ 50 0.4 2.275
+ 50 0.4 2.3
+ 50 0.4 2.325
+ 50 0.4 2.35
+ 50 0.4 2.375
+ 50 0.4 2.4
+ 50 0.4 2.425
+ 50 0.4 2.45
+ 50 0.4 2.475
+ 50 0.4 2.5
+ 52 0.4 1.25
+ 52 0.4 1.275
+ 52 0.4 1.3
+ 52 0.4 1.325
+ 52 0.4 1.35
+ 52 0.4 1.375
+ 52 0.4 1.4
+ 52 0.4 1.425
+ 52 0.4 1.45
+ 52 0.4 1.475
+ 52 0.4 1.5
+ 52 0.4 1.525
+ 52 0.4 1.55
+ 52 0.4 1.575
+ 52 0.4 1.6
+ 52 0.4 1.625
+ 52 0.4 1.65
+ 52 0.4 1.675
+ 52 0.4 1.7
+ 52 0.4 1.725
+ 52 0.4 1.75
+ 52 0.4 1.775
+ 52 0.4 1.8
+ 52 0.4 1.825
+ 52 0.4 1.85
+ 52 0.4 1.875
+ 52 0.4 1.9
+ 52 0.4 1.925
+ 52 0.4 1.95
+ 52 0.4 1.975
+ 52 0.4 2.0
+ 52 0.4 2.025
+ 52 0.4 2.05
+ 52 0.4 2.075
+ 52 0.4 2.1
+ 52 0.4 2.125
+ 52 0.4 2.15
+ 52 0.4 2.175
+ 52 0.4 2.2
+ 52 0.4 2.225
+ 52 0.4 2.25
+ 52 0.4 2.275
+ 52 0.4 2.3
+ 52 0.4 2.325
+ 52 0.4 2.35
+ 52 0.4 2.375
+ 52 0.4 2.4
+ 52 0.4 2.425
+ 52 0.4 2.45
+ 52 0.4 2.475
+ 52 0.4 2.5
+ 54 0.4 1.25
+ 54 0.4 1.275
+ 54 0.4 1.3
+ 54 0.4 1.325
+ 54 0.4 1.35
+ 54 0.4 1.375
+ 54 0.4 1.4
+ 54 0.4 1.425
+ 54 0.4 1.45
+ 54 0.4 1.475
+ 54 0.4 1.5
+ 54 0.4 1.525
+ 54 0.4 1.55
+ 54 0.4 1.575
+ 54 0.4 1.6
+ 54 0.4 1.625
+ 54 0.4 1.65
+ 54 0.4 1.675
+ 54 0.4 1.7
+ 54 0.4 1.725
+ 54 0.4 1.75
+ 54 0.4 1.775
+ 54 0.4 1.8
+ 54 0.4 1.825
+ 54 0.4 1.85
+ 54 0.4 1.875
+ 54 0.4 1.9
+ 54 0.4 1.925
+ 54 0.4 1.95
+ 54 0.4 1.975
+ 54 0.4 2.0
+ 54 0.4 2.025
+ 54 0.4 2.05
+ 54 0.4 2.075
+ 54 0.4 2.1
+ 54 0.4 2.125
+ 54 0.4 2.15
+ 54 0.4 2.175
+ 54 0.4 2.2
+ 54 0.4 2.225
+ 54 0.4 2.25
+ 54 0.4 2.275
+ 54 0.4 2.3
+ 54 0.4 2.325
+ 54 0.4 2.35
+ 54 0.4 2.375
+ 54 0.4 2.4
+ 54 0.4 2.425
+ 54 0.4 2.45
+ 54 0.4 2.475
+ 54 0.4 2.5
+ 56 0.4 1.25
+ 56 0.4 1.275
+ 56 0.4 1.3
+ 56 0.4 1.325
+ 56 0.4 1.35
+ 56 0.4 1.375
+ 56 0.4 1.4
+ 56 0.4 1.425
+ 56 0.4 1.45
+ 56 0.4 1.475
+ 56 0.4 1.5
+ 56 0.4 1.525
+ 56 0.4 1.55
+ 56 0.4 1.575
+ 56 0.4 1.6
+ 56 0.4 1.625
+ 56 0.4 1.65
+ 56 0.4 1.675
+ 56 0.4 1.7
+ 56 0.4 1.725
+ 56 0.4 1.75
+ 56 0.4 1.775
+ 56 0.4 1.8
+ 56 0.4 1.825
+ 56 0.4 1.85
+ 56 0.4 1.875
+ 56 0.4 1.9
+ 56 0.4 1.925
+ 56 0.4 1.95
+ 56 0.4 1.975
+ 56 0.4 2.0
+ 56 0.4 2.025
+ 56 0.4 2.05
+ 56 0.4 2.075
+ 56 0.4 2.1
+ 56 0.4 2.125
+ 56 0.4 2.15
+ 56 0.4 2.175
+ 56 0.4 2.2
+ 56 0.4 2.225
+ 56 0.4 2.25
+ 56 0.4 2.275
+ 56 0.4 2.3
+ 56 0.4 2.325
+ 56 0.4 2.35
+ 56 0.4 2.375
+ 56 0.4 2.4
+ 56 0.4 2.425
+ 56 0.4 2.45
+ 56 0.4 2.475
+ 56 0.4 2.5
+ 58 0.4 1.25
+ 58 0.4 1.275
+ 58 0.4 1.3
+ 58 0.4 1.325
+ 58 0.4 1.35
+ 58 0.4 1.375
+ 58 0.4 1.4
+ 58 0.4 1.425
+ 58 0.4 1.45
+ 58 0.4 1.475
+ 58 0.4 1.5
+ 58 0.4 1.525
+ 58 0.4 1.55
+ 58 0.4 1.575
+ 58 0.4 1.6
+ 58 0.4 1.625
+ 58 0.4 1.65
+ 58 0.4 1.675
+ 58 0.4 1.7
+ 58 0.4 1.725
+ 58 0.4 1.75
+ 58 0.4 1.775
+ 58 0.4 1.8
+ 58 0.4 1.825
+ 58 0.4 1.85
+ 58 0.4 1.875
+ 58 0.4 1.9
+ 58 0.4 1.925
+ 58 0.4 1.95
+ 58 0.4 1.975
+ 58 0.4 2.0
+ 58 0.4 2.025
+ 58 0.4 2.05
+ 58 0.4 2.075
+ 58 0.4 2.1
+ 58 0.4 2.125
+ 58 0.4 2.15
+ 58 0.4 2.175
+ 58 0.4 2.2
+ 58 0.4 2.225
+ 58 0.4 2.25
+ 58 0.4 2.275
+ 58 0.4 2.3
+ 58 0.4 2.325
+ 58 0.4 2.35
+ 58 0.4 2.375
+ 58 0.4 2.4
+ 58 0.4 2.425
+ 58 0.4 2.45
+ 58 0.4 2.475
+ 58 0.4 2.5
+ 60 0.4 1.25
+ 60 0.4 1.275
+ 60 0.4 1.3
+ 60 0.4 1.325
+ 60 0.4 1.35
+ 60 0.4 1.375
+ 60 0.4 1.4
+ 60 0.4 1.425
+ 60 0.4 1.45
+ 60 0.4 1.475
+ 60 0.4 1.5
+ 60 0.4 1.525
+ 60 0.4 1.55
+ 60 0.4 1.575
+ 60 0.4 1.6
+ 60 0.4 1.625
+ 60 0.4 1.65
+ 60 0.4 1.675
+ 60 0.4 1.7
+ 60 0.4 1.725
+ 60 0.4 1.75
+ 60 0.4 1.775
+ 60 0.4 1.8
+ 60 0.4 1.825
+ 60 0.4 1.85
+ 60 0.4 1.875
+ 60 0.4 1.9
+ 60 0.4 1.925
+ 60 0.4 1.95
+ 60 0.4 1.975
+ 60 0.4 2.0
+ 60 0.4 2.025
+ 60 0.4 2.05
+ 60 0.4 2.075
+ 60 0.4 2.1
+ 60 0.4 2.125
+ 60 0.4 2.15
+ 60 0.4 2.175
+ 60 0.4 2.2
+ 60 0.4 2.225
+ 60 0.4 2.25
+ 60 0.4 2.275
+ 60 0.4 2.3
+ 60 0.4 2.325
+ 60 0.4 2.35
+ 60 0.4 2.375
+ 60 0.4 2.4
+ 60 0.4 2.425
+ 60 0.4 2.45
+ 60 0.4 2.475
+ 60 0.4 2.5
+ 62 0.4 1.25
+ 62 0.4 1.275
+ 62 0.4 1.3
+ 62 0.4 1.325
+ 62 0.4 1.35
+ 62 0.4 1.375
+ 62 0.4 1.4
+ 62 0.4 1.425
+ 62 0.4 1.45
+ 62 0.4 1.475
+ 62 0.4 1.5
+ 62 0.4 1.525
+ 62 0.4 1.55
+ 62 0.4 1.575
+ 62 0.4 1.6
+ 62 0.4 1.625
+ 62 0.4 1.65
+ 62 0.4 1.675
+ 62 0.4 1.7
+ 62 0.4 1.725
+ 62 0.4 1.75
+ 62 0.4 1.775
+ 62 0.4 1.8
+ 62 0.4 1.825
+ 62 0.4 1.85
+ 62 0.4 1.875
+ 62 0.4 1.9
+ 62 0.4 1.925
+ 62 0.4 1.95
+ 62 0.4 1.975
+ 62 0.4 2.0
+ 62 0.4 2.025
+ 62 0.4 2.05
+ 62 0.4 2.075
+ 62 0.4 2.1
+ 62 0.4 2.125
+ 62 0.4 2.15
+ 62 0.4 2.175
+ 62 0.4 2.2
+ 62 0.4 2.225
+ 62 0.4 2.25
+ 62 0.4 2.275
+ 62 0.4 2.3
+ 62 0.4 2.325
+ 62 0.4 2.35
+ 62 0.4 2.375
+ 62 0.4 2.4
+ 62 0.4 2.425
+ 62 0.4 2.45
+ 62 0.4 2.475
+ 62 0.4 2.5
+ 64 0.4 1.25
+ 64 0.4 1.275
+ 64 0.4 1.3
+ 64 0.4 1.325
+ 64 0.4 1.35
+ 64 0.4 1.375
+ 64 0.4 1.4
+ 64 0.4 1.425
+ 64 0.4 1.45
+ 64 0.4 1.475
+ 64 0.4 1.5
+ 64 0.4 1.525
+ 64 0.4 1.55
+ 64 0.4 1.575
+ 64 0.4 1.6
+ 64 0.4 1.625
+ 64 0.4 1.65
+ 64 0.4 1.675
+ 64 0.4 1.7
+ 64 0.4 1.725
+ 64 0.4 1.75
+ 64 0.4 1.775
+ 64 0.4 1.8
+ 64 0.4 1.825
+ 64 0.4 1.85
+ 64 0.4 1.875
+ 64 0.4 1.9
+ 64 0.4 1.925
+ 64 0.4 1.95
+ 64 0.4 1.975
+ 64 0.4 2.0
+ 64 0.4 2.025
+ 64 0.4 2.05
+ 64 0.4 2.075
+ 64 0.4 2.1
+ 64 0.4 2.125
+ 64 0.4 2.15
+ 64 0.4 2.175
+ 64 0.4 2.2
+ 64 0.4 2.225
+ 64 0.4 2.25
+ 64 0.4 2.275
+ 64 0.4 2.3
+ 64 0.4 2.325
+ 64 0.4 2.35
+ 64 0.4 2.375
+ 64 0.4 2.4
+ 64 0.4 2.425
+ 64 0.4 2.45
+ 64 0.4 2.475
+ 64 0.4 2.5
+ 66 0.4 1.25
+ 66 0.4 1.275
+ 66 0.4 1.3
+ 66 0.4 1.325
+ 66 0.4 1.35
+ 66 0.4 1.375
+ 66 0.4 1.4
+ 66 0.4 1.425
+ 66 0.4 1.45
+ 66 0.4 1.475
+ 66 0.4 1.5
+ 66 0.4 1.525
+ 66 0.4 1.55
+ 66 0.4 1.575
+ 66 0.4 1.6
+ 66 0.4 1.625
+ 66 0.4 1.65
+ 66 0.4 1.675
+ 66 0.4 1.7
+ 66 0.4 1.725
+ 66 0.4 1.75
+ 66 0.4 1.775
+ 66 0.4 1.8
+ 66 0.4 1.825
+ 66 0.4 1.85
+ 66 0.4 1.875
+ 66 0.4 1.9
+ 66 0.4 1.925
+ 66 0.4 1.95
+ 66 0.4 1.975
+ 66 0.4 2.0
+ 66 0.4 2.025
+ 66 0.4 2.05
+ 66 0.4 2.075
+ 66 0.4 2.1
+ 66 0.4 2.125
+ 66 0.4 2.15
+ 66 0.4 2.175
+ 66 0.4 2.2
+ 66 0.4 2.225
+ 66 0.4 2.25
+ 66 0.4 2.275
+ 66 0.4 2.3
+ 66 0.4 2.325
+ 66 0.4 2.35
+ 66 0.4 2.375
+ 66 0.4 2.4
+ 66 0.4 2.425
+ 66 0.4 2.45
+ 66 0.4 2.475
+ 66 0.4 2.5
+ 68 0.4 1.25
+ 68 0.4 1.275
+ 68 0.4 1.3
+ 68 0.4 1.325
+ 68 0.4 1.35
+ 68 0.4 1.375
+ 68 0.4 1.4
+ 68 0.4 1.425
+ 68 0.4 1.45
+ 68 0.4 1.475
+ 68 0.4 1.5
+ 68 0.4 1.525
+ 68 0.4 1.55
+ 68 0.4 1.575
+ 68 0.4 1.6
+ 68 0.4 1.625
+ 68 0.4 1.65
+ 68 0.4 1.675
+ 68 0.4 1.7
+ 68 0.4 1.725
+ 68 0.4 1.75
+ 68 0.4 1.775
+ 68 0.4 1.8
+ 68 0.4 1.825
+ 68 0.4 1.85
+ 68 0.4 1.875
+ 68 0.4 1.9
+ 68 0.4 1.925
+ 68 0.4 1.95
+ 68 0.4 1.975
+ 68 0.4 2.0
+ 68 0.4 2.025
+ 68 0.4 2.05
+ 68 0.4 2.075
+ 68 0.4 2.1
+ 68 0.4 2.125
+ 68 0.4 2.15
+ 68 0.4 2.175
+ 68 0.4 2.2
+ 68 0.4 2.225
+ 68 0.4 2.25
+ 68 0.4 2.275
+ 68 0.4 2.3
+ 68 0.4 2.325
+ 68 0.4 2.35
+ 68 0.4 2.375
+ 68 0.4 2.4
+ 68 0.4 2.425
+ 68 0.4 2.45
+ 68 0.4 2.475
+ 68 0.4 2.5
+ 70 0.4 1.25
+ 70 0.4 1.275
+ 70 0.4 1.3
+ 70 0.4 1.325
+ 70 0.4 1.35
+ 70 0.4 1.375
+ 70 0.4 1.4
+ 70 0.4 1.425
+ 70 0.4 1.45
+ 70 0.4 1.475
+ 70 0.4 1.5
+ 70 0.4 1.525
+ 70 0.4 1.55
+ 70 0.4 1.575
+ 70 0.4 1.6
+ 70 0.4 1.625
+ 70 0.4 1.65
+ 70 0.4 1.675
+ 70 0.4 1.7
+ 70 0.4 1.725
+ 70 0.4 1.75
+ 70 0.4 1.775
+ 70 0.4 1.8
+ 70 0.4 1.825
+ 70 0.4 1.85
+ 70 0.4 1.875
+ 70 0.4 1.9
+ 70 0.4 1.925
+ 70 0.4 1.95
+ 70 0.4 1.975
+ 70 0.4 2.0
+ 70 0.4 2.025
+ 70 0.4 2.05
+ 70 0.4 2.075
+ 70 0.4 2.1
+ 70 0.4 2.125
+ 70 0.4 2.15
+ 70 0.4 2.175
+ 70 0.4 2.2
+ 70 0.4 2.225
+ 70 0.4 2.25
+ 70 0.4 2.275
+ 70 0.4 2.3
+ 70 0.4 2.325
+ 70 0.4 2.35
+ 70 0.4 2.375
+ 70 0.4 2.4
+ 70 0.4 2.425
+ 70 0.4 2.45
+ 70 0.4 2.475
+ 70 0.4 2.5
+ 72 0.4 1.25
+ 72 0.4 1.275
+ 72 0.4 1.3
+ 72 0.4 1.325
+ 72 0.4 1.35
+ 72 0.4 1.375
+ 72 0.4 1.4
+ 72 0.4 1.425
+ 72 0.4 1.45
+ 72 0.4 1.475
+ 72 0.4 1.5
+ 72 0.4 1.525
+ 72 0.4 1.55
+ 72 0.4 1.575
+ 72 0.4 1.6
+ 72 0.4 1.625
+ 72 0.4 1.65
+ 72 0.4 1.675
+ 72 0.4 1.7
+ 72 0.4 1.725
+ 72 0.4 1.75
+ 72 0.4 1.775
+ 72 0.4 1.8
+ 72 0.4 1.825
+ 72 0.4 1.85
+ 72 0.4 1.875
+ 72 0.4 1.9
+ 72 0.4 1.925
+ 72 0.4 1.95
+ 72 0.4 1.975
+ 72 0.4 2.0
+ 72 0.4 2.025
+ 72 0.4 2.05
+ 72 0.4 2.075
+ 72 0.4 2.1
+ 72 0.4 2.125
+ 72 0.4 2.15
+ 72 0.4 2.175
+ 72 0.4 2.2
+ 72 0.4 2.225
+ 72 0.4 2.25
+ 72 0.4 2.275
+ 72 0.4 2.3
+ 72 0.4 2.325
+ 72 0.4 2.35
+ 72 0.4 2.375
+ 72 0.4 2.4
+ 72 0.4 2.425
+ 72 0.4 2.45
+ 72 0.4 2.475
+ 72 0.4 2.5
+ 74 0.4 1.25
+ 74 0.4 1.275
+ 74 0.4 1.3
+ 74 0.4 1.325
+ 74 0.4 1.35
+ 74 0.4 1.375
+ 74 0.4 1.4
+ 74 0.4 1.425
+ 74 0.4 1.45
+ 74 0.4 1.475
+ 74 0.4 1.5
+ 74 0.4 1.525
+ 74 0.4 1.55
+ 74 0.4 1.575
+ 74 0.4 1.6
+ 74 0.4 1.625
+ 74 0.4 1.65
+ 74 0.4 1.675
+ 74 0.4 1.7
+ 74 0.4 1.725
+ 74 0.4 1.75
+ 74 0.4 1.775
+ 74 0.4 1.8
+ 74 0.4 1.825
+ 74 0.4 1.85
+ 74 0.4 1.875
+ 74 0.4 1.9
+ 74 0.4 1.925
+ 74 0.4 1.95
+ 74 0.4 1.975
+ 74 0.4 2.0
+ 74 0.4 2.025
+ 74 0.4 2.05
+ 74 0.4 2.075
+ 74 0.4 2.1
+ 74 0.4 2.125
+ 74 0.4 2.15
+ 74 0.4 2.175
+ 74 0.4 2.2
+ 74 0.4 2.225
+ 74 0.4 2.25
+ 74 0.4 2.275
+ 74 0.4 2.3
+ 74 0.4 2.325
+ 74 0.4 2.35
+ 74 0.4 2.375
+ 74 0.4 2.4
+ 74 0.4 2.425
+ 74 0.4 2.45
+ 74 0.4 2.475
+ 74 0.4 2.5
+ 76 0.4 1.25
+ 76 0.4 1.275
+ 76 0.4 1.3
+ 76 0.4 1.325
+ 76 0.4 1.35
+ 76 0.4 1.375
+ 76 0.4 1.4
+ 76 0.4 1.425
+ 76 0.4 1.45
+ 76 0.4 1.475
+ 76 0.4 1.5
+ 76 0.4 1.525
+ 76 0.4 1.55
+ 76 0.4 1.575
+ 76 0.4 1.6
+ 76 0.4 1.625
+ 76 0.4 1.65
+ 76 0.4 1.675
+ 76 0.4 1.7
+ 76 0.4 1.725
+ 76 0.4 1.75
+ 76 0.4 1.775
+ 76 0.4 1.8
+ 76 0.4 1.825
+ 76 0.4 1.85
+ 76 0.4 1.875
+ 76 0.4 1.9
+ 76 0.4 1.925
+ 76 0.4 1.95
+ 76 0.4 1.975
+ 76 0.4 2.0
+ 76 0.4 2.025
+ 76 0.4 2.05
+ 76 0.4 2.075
+ 76 0.4 2.1
+ 76 0.4 2.125
+ 76 0.4 2.15
+ 76 0.4 2.175
+ 76 0.4 2.2
+ 76 0.4 2.225
+ 76 0.4 2.25
+ 76 0.4 2.275
+ 76 0.4 2.3
+ 76 0.4 2.325
+ 76 0.4 2.35
+ 76 0.4 2.375
+ 76 0.4 2.4
+ 76 0.4 2.425
+ 76 0.4 2.45
+ 76 0.4 2.475
+ 76 0.4 2.5
+ 78 0.4 1.25
+ 78 0.4 1.275
+ 78 0.4 1.3
+ 78 0.4 1.325
+ 78 0.4 1.35
+ 78 0.4 1.375
+ 78 0.4 1.4
+ 78 0.4 1.425
+ 78 0.4 1.45
+ 78 0.4 1.475
+ 78 0.4 1.5
+ 78 0.4 1.525
+ 78 0.4 1.55
+ 78 0.4 1.575
+ 78 0.4 1.6
+ 78 0.4 1.625
+ 78 0.4 1.65
+ 78 0.4 1.675
+ 78 0.4 1.7
+ 78 0.4 1.725
+ 78 0.4 1.75
+ 78 0.4 1.775
+ 78 0.4 1.8
+ 78 0.4 1.825
+ 78 0.4 1.85
+ 78 0.4 1.875
+ 78 0.4 1.9
+ 78 0.4 1.925
+ 78 0.4 1.95
+ 78 0.4 1.975
+ 78 0.4 2.0
+ 78 0.4 2.025
+ 78 0.4 2.05
+ 78 0.4 2.075
+ 78 0.4 2.1
+ 78 0.4 2.125
+ 78 0.4 2.15
+ 78 0.4 2.175
+ 78 0.4 2.2
+ 78 0.4 2.225
+ 78 0.4 2.25
+ 78 0.4 2.275
+ 78 0.4 2.3
+ 78 0.4 2.325
+ 78 0.4 2.35
+ 78 0.4 2.375
+ 78 0.4 2.4
+ 78 0.4 2.425
+ 78 0.4 2.45
+ 78 0.4 2.475
+ 78 0.4 2.5
+ 80 0.4 1.25
+ 80 0.4 1.275
+ 80 0.4 1.3
+ 80 0.4 1.325
+ 80 0.4 1.35
+ 80 0.4 1.375
+ 80 0.4 1.4
+ 80 0.4 1.425
+ 80 0.4 1.45
+ 80 0.4 1.475
+ 80 0.4 1.5
+ 80 0.4 1.525
+ 80 0.4 1.55
+ 80 0.4 1.575
+ 80 0.4 1.6
+ 80 0.4 1.625
+ 80 0.4 1.65
+ 80 0.4 1.675
+ 80 0.4 1.7
+ 80 0.4 1.725
+ 80 0.4 1.75
+ 80 0.4 1.775
+ 80 0.4 1.8
+ 80 0.4 1.825
+ 80 0.4 1.85
+ 80 0.4 1.875
+ 80 0.4 1.9
+ 80 0.4 1.925
+ 80 0.4 1.95
+ 80 0.4 1.975
+ 80 0.4 2.0
+ 80 0.4 2.025
+ 80 0.4 2.05
+ 80 0.4 2.075
+ 80 0.4 2.1
+ 80 0.4 2.125
+ 80 0.4 2.15
+ 80 0.4 2.175
+ 80 0.4 2.2
+ 80 0.4 2.225
+ 80 0.4 2.25
+ 80 0.4 2.275
+ 80 0.4 2.3
+ 80 0.4 2.325
+ 80 0.4 2.35
+ 80 0.4 2.375
+ 80 0.4 2.4
+ 80 0.4 2.425
+ 80 0.4 2.45
+ 80 0.4 2.475
+ 80 0.4 2.5
+ 82 0.4 1.25
+ 82 0.4 1.275
+ 82 0.4 1.3
+ 82 0.4 1.325
+ 82 0.4 1.35
+ 82 0.4 1.375
+ 82 0.4 1.4
+ 82 0.4 1.425
+ 82 0.4 1.45
+ 82 0.4 1.475
+ 82 0.4 1.5
+ 82 0.4 1.525
+ 82 0.4 1.55
+ 82 0.4 1.575
+ 82 0.4 1.6
+ 82 0.4 1.625
+ 82 0.4 1.65
+ 82 0.4 1.675
+ 82 0.4 1.7
+ 82 0.4 1.725
+ 82 0.4 1.75
+ 82 0.4 1.775
+ 82 0.4 1.8
+ 82 0.4 1.825
+ 82 0.4 1.85
+ 82 0.4 1.875
+ 82 0.4 1.9
+ 82 0.4 1.925
+ 82 0.4 1.95
+ 82 0.4 1.975
+ 82 0.4 2.0
+ 82 0.4 2.025
+ 82 0.4 2.05
+ 82 0.4 2.075
+ 82 0.4 2.1
+ 82 0.4 2.125
+ 82 0.4 2.15
+ 82 0.4 2.175
+ 82 0.4 2.2
+ 82 0.4 2.225
+ 82 0.4 2.25
+ 82 0.4 2.275
+ 82 0.4 2.3
+ 82 0.4 2.325
+ 82 0.4 2.35
+ 82 0.4 2.375
+ 82 0.4 2.4
+ 82 0.4 2.425
+ 82 0.4 2.45
+ 82 0.4 2.475
+ 82 0.4 2.5
+ 84 0.4 1.25
+ 84 0.4 1.275
+ 84 0.4 1.3
+ 84 0.4 1.325
+ 84 0.4 1.35
+ 84 0.4 1.375
+ 84 0.4 1.4
+ 84 0.4 1.425
+ 84 0.4 1.45
+ 84 0.4 1.475
+ 84 0.4 1.5
+ 84 0.4 1.525
+ 84 0.4 1.55
+ 84 0.4 1.575
+ 84 0.4 1.6
+ 84 0.4 1.625
+ 84 0.4 1.65
+ 84 0.4 1.675
+ 84 0.4 1.7
+ 84 0.4 1.725
+ 84 0.4 1.75
+ 84 0.4 1.775
+ 84 0.4 1.8
+ 84 0.4 1.825
+ 84 0.4 1.85
+ 84 0.4 1.875
+ 84 0.4 1.9
+ 84 0.4 1.925
+ 84 0.4 1.95
+ 84 0.4 1.975
+ 84 0.4 2.0
+ 84 0.4 2.025
+ 84 0.4 2.05
+ 84 0.4 2.075
+ 84 0.4 2.1
+ 84 0.4 2.125
+ 84 0.4 2.15
+ 84 0.4 2.175
+ 84 0.4 2.2
+ 84 0.4 2.225
+ 84 0.4 2.25
+ 84 0.4 2.275
+ 84 0.4 2.3
+ 84 0.4 2.325
+ 84 0.4 2.35
+ 84 0.4 2.375
+ 84 0.4 2.4
+ 84 0.4 2.425
+ 84 0.4 2.45
+ 84 0.4 2.475
+ 84 0.4 2.5
+ 86 0.4 1.25
+ 86 0.4 1.275
+ 86 0.4 1.3
+ 86 0.4 1.325
+ 86 0.4 1.35
+ 86 0.4 1.375
+ 86 0.4 1.4
+ 86 0.4 1.425
+ 86 0.4 1.45
+ 86 0.4 1.475
+ 86 0.4 1.5
+ 86 0.4 1.525
+ 86 0.4 1.55
+ 86 0.4 1.575
+ 86 0.4 1.6
+ 86 0.4 1.625
+ 86 0.4 1.65
+ 86 0.4 1.675
+ 86 0.4 1.7
+ 86 0.4 1.725
+ 86 0.4 1.75
+ 86 0.4 1.775
+ 86 0.4 1.8
+ 86 0.4 1.825
+ 86 0.4 1.85
+ 86 0.4 1.875
+ 86 0.4 1.9
+ 86 0.4 1.925
+ 86 0.4 1.95
+ 86 0.4 1.975
+ 86 0.4 2.0
+ 86 0.4 2.025
+ 86 0.4 2.05
+ 86 0.4 2.075
+ 86 0.4 2.1
+ 86 0.4 2.125
+ 86 0.4 2.15
+ 86 0.4 2.175
+ 86 0.4 2.2
+ 86 0.4 2.225
+ 86 0.4 2.25
+ 86 0.4 2.275
+ 86 0.4 2.3
+ 86 0.4 2.325
+ 86 0.4 2.35
+ 86 0.4 2.375
+ 86 0.4 2.4
+ 86 0.4 2.425
+ 86 0.4 2.45
+ 86 0.4 2.475
+ 86 0.4 2.5
+ 88 0.4 1.25
+ 88 0.4 1.275
+ 88 0.4 1.3
+ 88 0.4 1.325
+ 88 0.4 1.35
+ 88 0.4 1.375
+ 88 0.4 1.4
+ 88 0.4 1.425
+ 88 0.4 1.45
+ 88 0.4 1.475
+ 88 0.4 1.5
+ 88 0.4 1.525
+ 88 0.4 1.55
+ 88 0.4 1.575
+ 88 0.4 1.6
+ 88 0.4 1.625
+ 88 0.4 1.65
+ 88 0.4 1.675
+ 88 0.4 1.7
+ 88 0.4 1.725
+ 88 0.4 1.75
+ 88 0.4 1.775
+ 88 0.4 1.8
+ 88 0.4 1.825
+ 88 0.4 1.85
+ 88 0.4 1.875
+ 88 0.4 1.9
+ 88 0.4 1.925
+ 88 0.4 1.95
+ 88 0.4 1.975
+ 88 0.4 2.0
+ 88 0.4 2.025
+ 88 0.4 2.05
+ 88 0.4 2.075
+ 88 0.4 2.1
+ 88 0.4 2.125
+ 88 0.4 2.15
+ 88 0.4 2.175
+ 88 0.4 2.2
+ 88 0.4 2.225
+ 88 0.4 2.25
+ 88 0.4 2.275
+ 88 0.4 2.3
+ 88 0.4 2.325
+ 88 0.4 2.35
+ 88 0.4 2.375
+ 88 0.4 2.4
+ 88 0.4 2.425
+ 88 0.4 2.45
+ 88 0.4 2.475
+ 88 0.4 2.5
+ 90 0.4 1.25
+ 90 0.4 1.275
+ 90 0.4 1.3
+ 90 0.4 1.325
+ 90 0.4 1.35
+ 90 0.4 1.375
+ 90 0.4 1.4
+ 90 0.4 1.425
+ 90 0.4 1.45
+ 90 0.4 1.475
+ 90 0.4 1.5
+ 90 0.4 1.525
+ 90 0.4 1.55
+ 90 0.4 1.575
+ 90 0.4 1.6
+ 90 0.4 1.625
+ 90 0.4 1.65
+ 90 0.4 1.675
+ 90 0.4 1.7
+ 90 0.4 1.725
+ 90 0.4 1.75
+ 90 0.4 1.775
+ 90 0.4 1.8
+ 90 0.4 1.825
+ 90 0.4 1.85
+ 90 0.4 1.875
+ 90 0.4 1.9
+ 90 0.4 1.925
+ 90 0.4 1.95
+ 90 0.4 1.975
+ 90 0.4 2.0
+ 90 0.4 2.025
+ 90 0.4 2.05
+ 90 0.4 2.075
+ 90 0.4 2.1
+ 90 0.4 2.125
+ 90 0.4 2.15
+ 90 0.4 2.175
+ 90 0.4 2.2
+ 90 0.4 2.225
+ 90 0.4 2.25
+ 90 0.4 2.275
+ 90 0.4 2.3
+ 90 0.4 2.325
+ 90 0.4 2.35
+ 90 0.4 2.375
+ 90 0.4 2.4
+ 90 0.4 2.425
+ 90 0.4 2.45
+ 90 0.4 2.475
+ 90 0.4 2.5
+ 92 0.4 1.25
+ 92 0.4 1.275
+ 92 0.4 1.3
+ 92 0.4 1.325
+ 92 0.4 1.35
+ 92 0.4 1.375
+ 92 0.4 1.4
+ 92 0.4 1.425
+ 92 0.4 1.45
+ 92 0.4 1.475
+ 92 0.4 1.5
+ 92 0.4 1.525
+ 92 0.4 1.55
+ 92 0.4 1.575
+ 92 0.4 1.6
+ 92 0.4 1.625
+ 92 0.4 1.65
+ 92 0.4 1.675
+ 92 0.4 1.7
+ 92 0.4 1.725
+ 92 0.4 1.75
+ 92 0.4 1.775
+ 92 0.4 1.8
+ 92 0.4 1.825
+ 92 0.4 1.85
+ 92 0.4 1.875
+ 92 0.4 1.9
+ 92 0.4 1.925
+ 92 0.4 1.95
+ 92 0.4 1.975
+ 92 0.4 2.0
+ 92 0.4 2.025
+ 92 0.4 2.05
+ 92 0.4 2.075
+ 92 0.4 2.1
+ 92 0.4 2.125
+ 92 0.4 2.15
+ 92 0.4 2.175
+ 92 0.4 2.2
+ 92 0.4 2.225
+ 92 0.4 2.25
+ 92 0.4 2.275
+ 92 0.4 2.3
+ 92 0.4 2.325
+ 92 0.4 2.35
+ 92 0.4 2.375
+ 92 0.4 2.4
+ 92 0.4 2.425
+ 92 0.4 2.45
+ 92 0.4 2.475
+ 92 0.4 2.5
+ 94 0.4 1.25
+ 94 0.4 1.275
+ 94 0.4 1.3
+ 94 0.4 1.325
+ 94 0.4 1.35
+ 94 0.4 1.375
+ 94 0.4 1.4
+ 94 0.4 1.425
+ 94 0.4 1.45
+ 94 0.4 1.475
+ 94 0.4 1.5
+ 94 0.4 1.525
+ 94 0.4 1.55
+ 94 0.4 1.575
+ 94 0.4 1.6
+ 94 0.4 1.625
+ 94 0.4 1.65
+ 94 0.4 1.675
+ 94 0.4 1.7
+ 94 0.4 1.725
+ 94 0.4 1.75
+ 94 0.4 1.775
+ 94 0.4 1.8
+ 94 0.4 1.825
+ 94 0.4 1.85
+ 94 0.4 1.875
+ 94 0.4 1.9
+ 94 0.4 1.925
+ 94 0.4 1.95
+ 94 0.4 1.975
+ 94 0.4 2.0
+ 94 0.4 2.025
+ 94 0.4 2.05
+ 94 0.4 2.075
+ 94 0.4 2.1
+ 94 0.4 2.125
+ 94 0.4 2.15
+ 94 0.4 2.175
+ 94 0.4 2.2
+ 94 0.4 2.225
+ 94 0.4 2.25
+ 94 0.4 2.275
+ 94 0.4 2.3
+ 94 0.4 2.325
+ 94 0.4 2.35
+ 94 0.4 2.375
+ 94 0.4 2.4
+ 94 0.4 2.425
+ 94 0.4 2.45
+ 94 0.4 2.475
+ 94 0.4 2.5
+ 96 0.4 1.25
+ 96 0.4 1.275
+ 96 0.4 1.3
+ 96 0.4 1.325
+ 96 0.4 1.35
+ 96 0.4 1.375
+ 96 0.4 1.4
+ 96 0.4 1.425
+ 96 0.4 1.45
+ 96 0.4 1.475
+ 96 0.4 1.5
+ 96 0.4 1.525
+ 96 0.4 1.55
+ 96 0.4 1.575
+ 96 0.4 1.6
+ 96 0.4 1.625
+ 96 0.4 1.65
+ 96 0.4 1.675
+ 96 0.4 1.7
+ 96 0.4 1.725
+ 96 0.4 1.75
+ 96 0.4 1.775
+ 96 0.4 1.8
+ 96 0.4 1.825
+ 96 0.4 1.85
+ 96 0.4 1.875
+ 96 0.4 1.9
+ 96 0.4 1.925
+ 96 0.4 1.95
+ 96 0.4 1.975
+ 96 0.4 2.0
+ 96 0.4 2.025
+ 96 0.4 2.05
+ 96 0.4 2.075
+ 96 0.4 2.1
+ 96 0.4 2.125
+ 96 0.4 2.15
+ 96 0.4 2.175
+ 96 0.4 2.2
+ 96 0.4 2.225
+ 96 0.4 2.25
+ 96 0.4 2.275
+ 96 0.4 2.3
+ 96 0.4 2.325
+ 96 0.4 2.35
+ 96 0.4 2.375
+ 96 0.4 2.4
+ 96 0.4 2.425
+ 96 0.4 2.45
+ 96 0.4 2.475
+ 96 0.4 2.5
+ 98 0.4 1.25
+ 98 0.4 1.275
+ 98 0.4 1.3
+ 98 0.4 1.325
+ 98 0.4 1.35
+ 98 0.4 1.375
+ 98 0.4 1.4
+ 98 0.4 1.425
+ 98 0.4 1.45
+ 98 0.4 1.475
+ 98 0.4 1.5
+ 98 0.4 1.525
+ 98 0.4 1.55
+ 98 0.4 1.575
+ 98 0.4 1.6
+ 98 0.4 1.625
+ 98 0.4 1.65
+ 98 0.4 1.675
+ 98 0.4 1.7
+ 98 0.4 1.725
+ 98 0.4 1.75
+ 98 0.4 1.775
+ 98 0.4 1.8
+ 98 0.4 1.825
+ 98 0.4 1.85
+ 98 0.4 1.875
+ 98 0.4 1.9
+ 98 0.4 1.925
+ 98 0.4 1.95
+ 98 0.4 1.975
+ 98 0.4 2.0
+ 98 0.4 2.025
+ 98 0.4 2.05
+ 98 0.4 2.075
+ 98 0.4 2.1
+ 98 0.4 2.125
+ 98 0.4 2.15
+ 98 0.4 2.175
+ 98 0.4 2.2
+ 98 0.4 2.225
+ 98 0.4 2.25
+ 98 0.4 2.275
+ 98 0.4 2.3
+ 98 0.4 2.325
+ 98 0.4 2.35
+ 98 0.4 2.375
+ 98 0.4 2.4
+ 98 0.4 2.425
+ 98 0.4 2.45
+ 98 0.4 2.475
+ 98 0.4 2.5
+ 100 0.4 1.25
+ 100 0.4 1.275
+ 100 0.4 1.3
+ 100 0.4 1.325
+ 100 0.4 1.35
+ 100 0.4 1.375
+ 100 0.4 1.4
+ 100 0.4 1.425
+ 100 0.4 1.45
+ 100 0.4 1.475
+ 100 0.4 1.5
+ 100 0.4 1.525
+ 100 0.4 1.55
+ 100 0.4 1.575
+ 100 0.4 1.6
+ 100 0.4 1.625
+ 100 0.4 1.65
+ 100 0.4 1.675
+ 100 0.4 1.7
+ 100 0.4 1.725
+ 100 0.4 1.75
+ 100 0.4 1.775
+ 100 0.4 1.8
+ 100 0.4 1.825
+ 100 0.4 1.85
+ 100 0.4 1.875
+ 100 0.4 1.9
+ 100 0.4 1.925
+ 100 0.4 1.95
+ 100 0.4 1.975
+ 100 0.4 2.0
+ 100 0.4 2.025
+ 100 0.4 2.05
+ 100 0.4 2.075
+ 100 0.4 2.1
+ 100 0.4 2.125
+ 100 0.4 2.15
+ 100 0.4 2.175
+ 100 0.4 2.2
+ 100 0.4 2.225
+ 100 0.4 2.25
+ 100 0.4 2.275
+ 100 0.4 2.3
+ 100 0.4 2.325
+ 100 0.4 2.35
+ 100 0.4 2.375
+ 100 0.4 2.4
+ 100 0.4 2.425
+ 100 0.4 2.45
+ 100 0.4 2.475
+ 100 0.4 2.5
+ 0 0.5 1.25
+ 0 0.5 1.275
+ 0 0.5 1.3
+ 0 0.5 1.325
+ 0 0.5 1.35
+ 0 0.5 1.375
+ 0 0.5 1.4
+ 0 0.5 1.425
+ 0 0.5 1.45
+ 0 0.5 1.475
+ 0 0.5 1.5
+ 0 0.5 1.525
+ 0 0.5 1.55
+ 0 0.5 1.575
+ 0 0.5 1.6
+ 0 0.5 1.625
+ 0 0.5 1.65
+ 0 0.5 1.675
+ 0 0.5 1.7
+ 0 0.5 1.725
+ 0 0.5 1.75
+ 0 0.5 1.775
+ 0 0.5 1.8
+ 0 0.5 1.825
+ 0 0.5 1.85
+ 0 0.5 1.875
+ 0 0.5 1.9
+ 0 0.5 1.925
+ 0 0.5 1.95
+ 0 0.5 1.975
+ 0 0.5 2.0
+ 0 0.5 2.025
+ 0 0.5 2.05
+ 0 0.5 2.075
+ 0 0.5 2.1
+ 0 0.5 2.125
+ 0 0.5 2.15
+ 0 0.5 2.175
+ 0 0.5 2.2
+ 0 0.5 2.225
+ 0 0.5 2.25
+ 0 0.5 2.275
+ 0 0.5 2.3
+ 0 0.5 2.325
+ 0 0.5 2.35
+ 0 0.5 2.375
+ 0 0.5 2.4
+ 0 0.5 2.425
+ 0 0.5 2.45
+ 0 0.5 2.475
+ 0 0.5 2.5
+ 2 0.5 1.25
+ 2 0.5 1.275
+ 2 0.5 1.3
+ 2 0.5 1.325
+ 2 0.5 1.35
+ 2 0.5 1.375
+ 2 0.5 1.4
+ 2 0.5 1.425
+ 2 0.5 1.45
+ 2 0.5 1.475
+ 2 0.5 1.5
+ 2 0.5 1.525
+ 2 0.5 1.55
+ 2 0.5 1.575
+ 2 0.5 1.6
+ 2 0.5 1.625
+ 2 0.5 1.65
+ 2 0.5 1.675
+ 2 0.5 1.7
+ 2 0.5 1.725
+ 2 0.5 1.75
+ 2 0.5 1.775
+ 2 0.5 1.8
+ 2 0.5 1.825
+ 2 0.5 1.85
+ 2 0.5 1.875
+ 2 0.5 1.9
+ 2 0.5 1.925
+ 2 0.5 1.95
+ 2 0.5 1.975
+ 2 0.5 2.0
+ 2 0.5 2.025
+ 2 0.5 2.05
+ 2 0.5 2.075
+ 2 0.5 2.1
+ 2 0.5 2.125
+ 2 0.5 2.15
+ 2 0.5 2.175
+ 2 0.5 2.2
+ 2 0.5 2.225
+ 2 0.5 2.25
+ 2 0.5 2.275
+ 2 0.5 2.3
+ 2 0.5 2.325
+ 2 0.5 2.35
+ 2 0.5 2.375
+ 2 0.5 2.4
+ 2 0.5 2.425
+ 2 0.5 2.45
+ 2 0.5 2.475
+ 2 0.5 2.5
+ 4 0.5 1.25
+ 4 0.5 1.275
+ 4 0.5 1.3
+ 4 0.5 1.325
+ 4 0.5 1.35
+ 4 0.5 1.375
+ 4 0.5 1.4
+ 4 0.5 1.425
+ 4 0.5 1.45
+ 4 0.5 1.475
+ 4 0.5 1.5
+ 4 0.5 1.525
+ 4 0.5 1.55
+ 4 0.5 1.575
+ 4 0.5 1.6
+ 4 0.5 1.625
+ 4 0.5 1.65
+ 4 0.5 1.675
+ 4 0.5 1.7
+ 4 0.5 1.725
+ 4 0.5 1.75
+ 4 0.5 1.775
+ 4 0.5 1.8
+ 4 0.5 1.825
+ 4 0.5 1.85
+ 4 0.5 1.875
+ 4 0.5 1.9
+ 4 0.5 1.925
+ 4 0.5 1.95
+ 4 0.5 1.975
+ 4 0.5 2.0
+ 4 0.5 2.025
+ 4 0.5 2.05
+ 4 0.5 2.075
+ 4 0.5 2.1
+ 4 0.5 2.125
+ 4 0.5 2.15
+ 4 0.5 2.175
+ 4 0.5 2.2
+ 4 0.5 2.225
+ 4 0.5 2.25
+ 4 0.5 2.275
+ 4 0.5 2.3
+ 4 0.5 2.325
+ 4 0.5 2.35
+ 4 0.5 2.375
+ 4 0.5 2.4
+ 4 0.5 2.425
+ 4 0.5 2.45
+ 4 0.5 2.475
+ 4 0.5 2.5
+ 6 0.5 1.25
+ 6 0.5 1.275
+ 6 0.5 1.3
+ 6 0.5 1.325
+ 6 0.5 1.35
+ 6 0.5 1.375
+ 6 0.5 1.4
+ 6 0.5 1.425
+ 6 0.5 1.45
+ 6 0.5 1.475
+ 6 0.5 1.5
+ 6 0.5 1.525
+ 6 0.5 1.55
+ 6 0.5 1.575
+ 6 0.5 1.6
+ 6 0.5 1.625
+ 6 0.5 1.65
+ 6 0.5 1.675
+ 6 0.5 1.7
+ 6 0.5 1.725
+ 6 0.5 1.75
+ 6 0.5 1.775
+ 6 0.5 1.8
+ 6 0.5 1.825
+ 6 0.5 1.85
+ 6 0.5 1.875
+ 6 0.5 1.9
+ 6 0.5 1.925
+ 6 0.5 1.95
+ 6 0.5 1.975
+ 6 0.5 2.0
+ 6 0.5 2.025
+ 6 0.5 2.05
+ 6 0.5 2.075
+ 6 0.5 2.1
+ 6 0.5 2.125
+ 6 0.5 2.15
+ 6 0.5 2.175
+ 6 0.5 2.2
+ 6 0.5 2.225
+ 6 0.5 2.25
+ 6 0.5 2.275
+ 6 0.5 2.3
+ 6 0.5 2.325
+ 6 0.5 2.35
+ 6 0.5 2.375
+ 6 0.5 2.4
+ 6 0.5 2.425
+ 6 0.5 2.45
+ 6 0.5 2.475
+ 6 0.5 2.5
+ 8 0.5 1.25
+ 8 0.5 1.275
+ 8 0.5 1.3
+ 8 0.5 1.325
+ 8 0.5 1.35
+ 8 0.5 1.375
+ 8 0.5 1.4
+ 8 0.5 1.425
+ 8 0.5 1.45
+ 8 0.5 1.475
+ 8 0.5 1.5
+ 8 0.5 1.525
+ 8 0.5 1.55
+ 8 0.5 1.575
+ 8 0.5 1.6
+ 8 0.5 1.625
+ 8 0.5 1.65
+ 8 0.5 1.675
+ 8 0.5 1.7
+ 8 0.5 1.725
+ 8 0.5 1.75
+ 8 0.5 1.775
+ 8 0.5 1.8
+ 8 0.5 1.825
+ 8 0.5 1.85
+ 8 0.5 1.875
+ 8 0.5 1.9
+ 8 0.5 1.925
+ 8 0.5 1.95
+ 8 0.5 1.975
+ 8 0.5 2.0
+ 8 0.5 2.025
+ 8 0.5 2.05
+ 8 0.5 2.075
+ 8 0.5 2.1
+ 8 0.5 2.125
+ 8 0.5 2.15
+ 8 0.5 2.175
+ 8 0.5 2.2
+ 8 0.5 2.225
+ 8 0.5 2.25
+ 8 0.5 2.275
+ 8 0.5 2.3
+ 8 0.5 2.325
+ 8 0.5 2.35
+ 8 0.5 2.375
+ 8 0.5 2.4
+ 8 0.5 2.425
+ 8 0.5 2.45
+ 8 0.5 2.475
+ 8 0.5 2.5
+ 10 0.5 1.25
+ 10 0.5 1.275
+ 10 0.5 1.3
+ 10 0.5 1.325
+ 10 0.5 1.35
+ 10 0.5 1.375
+ 10 0.5 1.4
+ 10 0.5 1.425
+ 10 0.5 1.45
+ 10 0.5 1.475
+ 10 0.5 1.5
+ 10 0.5 1.525
+ 10 0.5 1.55
+ 10 0.5 1.575
+ 10 0.5 1.6
+ 10 0.5 1.625
+ 10 0.5 1.65
+ 10 0.5 1.675
+ 10 0.5 1.7
+ 10 0.5 1.725
+ 10 0.5 1.75
+ 10 0.5 1.775
+ 10 0.5 1.8
+ 10 0.5 1.825
+ 10 0.5 1.85
+ 10 0.5 1.875
+ 10 0.5 1.9
+ 10 0.5 1.925
+ 10 0.5 1.95
+ 10 0.5 1.975
+ 10 0.5 2.0
+ 10 0.5 2.025
+ 10 0.5 2.05
+ 10 0.5 2.075
+ 10 0.5 2.1
+ 10 0.5 2.125
+ 10 0.5 2.15
+ 10 0.5 2.175
+ 10 0.5 2.2
+ 10 0.5 2.225
+ 10 0.5 2.25
+ 10 0.5 2.275
+ 10 0.5 2.3
+ 10 0.5 2.325
+ 10 0.5 2.35
+ 10 0.5 2.375
+ 10 0.5 2.4
+ 10 0.5 2.425
+ 10 0.5 2.45
+ 10 0.5 2.475
+ 10 0.5 2.5
+ 12 0.5 1.25
+ 12 0.5 1.275
+ 12 0.5 1.3
+ 12 0.5 1.325
+ 12 0.5 1.35
+ 12 0.5 1.375
+ 12 0.5 1.4
+ 12 0.5 1.425
+ 12 0.5 1.45
+ 12 0.5 1.475
+ 12 0.5 1.5
+ 12 0.5 1.525
+ 12 0.5 1.55
+ 12 0.5 1.575
+ 12 0.5 1.6
+ 12 0.5 1.625
+ 12 0.5 1.65
+ 12 0.5 1.675
+ 12 0.5 1.7
+ 12 0.5 1.725
+ 12 0.5 1.75
+ 12 0.5 1.775
+ 12 0.5 1.8
+ 12 0.5 1.825
+ 12 0.5 1.85
+ 12 0.5 1.875
+ 12 0.5 1.9
+ 12 0.5 1.925
+ 12 0.5 1.95
+ 12 0.5 1.975
+ 12 0.5 2.0
+ 12 0.5 2.025
+ 12 0.5 2.05
+ 12 0.5 2.075
+ 12 0.5 2.1
+ 12 0.5 2.125
+ 12 0.5 2.15
+ 12 0.5 2.175
+ 12 0.5 2.2
+ 12 0.5 2.225
+ 12 0.5 2.25
+ 12 0.5 2.275
+ 12 0.5 2.3
+ 12 0.5 2.325
+ 12 0.5 2.35
+ 12 0.5 2.375
+ 12 0.5 2.4
+ 12 0.5 2.425
+ 12 0.5 2.45
+ 12 0.5 2.475
+ 12 0.5 2.5
+ 14 0.5 1.25
+ 14 0.5 1.275
+ 14 0.5 1.3
+ 14 0.5 1.325
+ 14 0.5 1.35
+ 14 0.5 1.375
+ 14 0.5 1.4
+ 14 0.5 1.425
+ 14 0.5 1.45
+ 14 0.5 1.475
+ 14 0.5 1.5
+ 14 0.5 1.525
+ 14 0.5 1.55
+ 14 0.5 1.575
+ 14 0.5 1.6
+ 14 0.5 1.625
+ 14 0.5 1.65
+ 14 0.5 1.675
+ 14 0.5 1.7
+ 14 0.5 1.725
+ 14 0.5 1.75
+ 14 0.5 1.775
+ 14 0.5 1.8
+ 14 0.5 1.825
+ 14 0.5 1.85
+ 14 0.5 1.875
+ 14 0.5 1.9
+ 14 0.5 1.925
+ 14 0.5 1.95
+ 14 0.5 1.975
+ 14 0.5 2.0
+ 14 0.5 2.025
+ 14 0.5 2.05
+ 14 0.5 2.075
+ 14 0.5 2.1
+ 14 0.5 2.125
+ 14 0.5 2.15
+ 14 0.5 2.175
+ 14 0.5 2.2
+ 14 0.5 2.225
+ 14 0.5 2.25
+ 14 0.5 2.275
+ 14 0.5 2.3
+ 14 0.5 2.325
+ 14 0.5 2.35
+ 14 0.5 2.375
+ 14 0.5 2.4
+ 14 0.5 2.425
+ 14 0.5 2.45
+ 14 0.5 2.475
+ 14 0.5 2.5
+ 16 0.5 1.25
+ 16 0.5 1.275
+ 16 0.5 1.3
+ 16 0.5 1.325
+ 16 0.5 1.35
+ 16 0.5 1.375
+ 16 0.5 1.4
+ 16 0.5 1.425
+ 16 0.5 1.45
+ 16 0.5 1.475
+ 16 0.5 1.5
+ 16 0.5 1.525
+ 16 0.5 1.55
+ 16 0.5 1.575
+ 16 0.5 1.6
+ 16 0.5 1.625
+ 16 0.5 1.65
+ 16 0.5 1.675
+ 16 0.5 1.7
+ 16 0.5 1.725
+ 16 0.5 1.75
+ 16 0.5 1.775
+ 16 0.5 1.8
+ 16 0.5 1.825
+ 16 0.5 1.85
+ 16 0.5 1.875
+ 16 0.5 1.9
+ 16 0.5 1.925
+ 16 0.5 1.95
+ 16 0.5 1.975
+ 16 0.5 2.0
+ 16 0.5 2.025
+ 16 0.5 2.05
+ 16 0.5 2.075
+ 16 0.5 2.1
+ 16 0.5 2.125
+ 16 0.5 2.15
+ 16 0.5 2.175
+ 16 0.5 2.2
+ 16 0.5 2.225
+ 16 0.5 2.25
+ 16 0.5 2.275
+ 16 0.5 2.3
+ 16 0.5 2.325
+ 16 0.5 2.35
+ 16 0.5 2.375
+ 16 0.5 2.4
+ 16 0.5 2.425
+ 16 0.5 2.45
+ 16 0.5 2.475
+ 16 0.5 2.5
+ 18 0.5 1.25
+ 18 0.5 1.275
+ 18 0.5 1.3
+ 18 0.5 1.325
+ 18 0.5 1.35
+ 18 0.5 1.375
+ 18 0.5 1.4
+ 18 0.5 1.425
+ 18 0.5 1.45
+ 18 0.5 1.475
+ 18 0.5 1.5
+ 18 0.5 1.525
+ 18 0.5 1.55
+ 18 0.5 1.575
+ 18 0.5 1.6
+ 18 0.5 1.625
+ 18 0.5 1.65
+ 18 0.5 1.675
+ 18 0.5 1.7
+ 18 0.5 1.725
+ 18 0.5 1.75
+ 18 0.5 1.775
+ 18 0.5 1.8
+ 18 0.5 1.825
+ 18 0.5 1.85
+ 18 0.5 1.875
+ 18 0.5 1.9
+ 18 0.5 1.925
+ 18 0.5 1.95
+ 18 0.5 1.975
+ 18 0.5 2.0
+ 18 0.5 2.025
+ 18 0.5 2.05
+ 18 0.5 2.075
+ 18 0.5 2.1
+ 18 0.5 2.125
+ 18 0.5 2.15
+ 18 0.5 2.175
+ 18 0.5 2.2
+ 18 0.5 2.225
+ 18 0.5 2.25
+ 18 0.5 2.275
+ 18 0.5 2.3
+ 18 0.5 2.325
+ 18 0.5 2.35
+ 18 0.5 2.375
+ 18 0.5 2.4
+ 18 0.5 2.425
+ 18 0.5 2.45
+ 18 0.5 2.475
+ 18 0.5 2.5
+ 20 0.5 1.25
+ 20 0.5 1.275
+ 20 0.5 1.3
+ 20 0.5 1.325
+ 20 0.5 1.35
+ 20 0.5 1.375
+ 20 0.5 1.4
+ 20 0.5 1.425
+ 20 0.5 1.45
+ 20 0.5 1.475
+ 20 0.5 1.5
+ 20 0.5 1.525
+ 20 0.5 1.55
+ 20 0.5 1.575
+ 20 0.5 1.6
+ 20 0.5 1.625
+ 20 0.5 1.65
+ 20 0.5 1.675
+ 20 0.5 1.7
+ 20 0.5 1.725
+ 20 0.5 1.75
+ 20 0.5 1.775
+ 20 0.5 1.8
+ 20 0.5 1.825
+ 20 0.5 1.85
+ 20 0.5 1.875
+ 20 0.5 1.9
+ 20 0.5 1.925
+ 20 0.5 1.95
+ 20 0.5 1.975
+ 20 0.5 2.0
+ 20 0.5 2.025
+ 20 0.5 2.05
+ 20 0.5 2.075
+ 20 0.5 2.1
+ 20 0.5 2.125
+ 20 0.5 2.15
+ 20 0.5 2.175
+ 20 0.5 2.2
+ 20 0.5 2.225
+ 20 0.5 2.25
+ 20 0.5 2.275
+ 20 0.5 2.3
+ 20 0.5 2.325
+ 20 0.5 2.35
+ 20 0.5 2.375
+ 20 0.5 2.4
+ 20 0.5 2.425
+ 20 0.5 2.45
+ 20 0.5 2.475
+ 20 0.5 2.5
+ 22 0.5 1.25
+ 22 0.5 1.275
+ 22 0.5 1.3
+ 22 0.5 1.325
+ 22 0.5 1.35
+ 22 0.5 1.375
+ 22 0.5 1.4
+ 22 0.5 1.425
+ 22 0.5 1.45
+ 22 0.5 1.475
+ 22 0.5 1.5
+ 22 0.5 1.525
+ 22 0.5 1.55
+ 22 0.5 1.575
+ 22 0.5 1.6
+ 22 0.5 1.625
+ 22 0.5 1.65
+ 22 0.5 1.675
+ 22 0.5 1.7
+ 22 0.5 1.725
+ 22 0.5 1.75
+ 22 0.5 1.775
+ 22 0.5 1.8
+ 22 0.5 1.825
+ 22 0.5 1.85
+ 22 0.5 1.875
+ 22 0.5 1.9
+ 22 0.5 1.925
+ 22 0.5 1.95
+ 22 0.5 1.975
+ 22 0.5 2.0
+ 22 0.5 2.025
+ 22 0.5 2.05
+ 22 0.5 2.075
+ 22 0.5 2.1
+ 22 0.5 2.125
+ 22 0.5 2.15
+ 22 0.5 2.175
+ 22 0.5 2.2
+ 22 0.5 2.225
+ 22 0.5 2.25
+ 22 0.5 2.275
+ 22 0.5 2.3
+ 22 0.5 2.325
+ 22 0.5 2.35
+ 22 0.5 2.375
+ 22 0.5 2.4
+ 22 0.5 2.425
+ 22 0.5 2.45
+ 22 0.5 2.475
+ 22 0.5 2.5
+ 24 0.5 1.25
+ 24 0.5 1.275
+ 24 0.5 1.3
+ 24 0.5 1.325
+ 24 0.5 1.35
+ 24 0.5 1.375
+ 24 0.5 1.4
+ 24 0.5 1.425
+ 24 0.5 1.45
+ 24 0.5 1.475
+ 24 0.5 1.5
+ 24 0.5 1.525
+ 24 0.5 1.55
+ 24 0.5 1.575
+ 24 0.5 1.6
+ 24 0.5 1.625
+ 24 0.5 1.65
+ 24 0.5 1.675
+ 24 0.5 1.7
+ 24 0.5 1.725
+ 24 0.5 1.75
+ 24 0.5 1.775
+ 24 0.5 1.8
+ 24 0.5 1.825
+ 24 0.5 1.85
+ 24 0.5 1.875
+ 24 0.5 1.9
+ 24 0.5 1.925
+ 24 0.5 1.95
+ 24 0.5 1.975
+ 24 0.5 2.0
+ 24 0.5 2.025
+ 24 0.5 2.05
+ 24 0.5 2.075
+ 24 0.5 2.1
+ 24 0.5 2.125
+ 24 0.5 2.15
+ 24 0.5 2.175
+ 24 0.5 2.2
+ 24 0.5 2.225
+ 24 0.5 2.25
+ 24 0.5 2.275
+ 24 0.5 2.3
+ 24 0.5 2.325
+ 24 0.5 2.35
+ 24 0.5 2.375
+ 24 0.5 2.4
+ 24 0.5 2.425
+ 24 0.5 2.45
+ 24 0.5 2.475
+ 24 0.5 2.5
+ 26 0.5 1.25
+ 26 0.5 1.275
+ 26 0.5 1.3
+ 26 0.5 1.325
+ 26 0.5 1.35
+ 26 0.5 1.375
+ 26 0.5 1.4
+ 26 0.5 1.425
+ 26 0.5 1.45
+ 26 0.5 1.475
+ 26 0.5 1.5
+ 26 0.5 1.525
+ 26 0.5 1.55
+ 26 0.5 1.575
+ 26 0.5 1.6
+ 26 0.5 1.625
+ 26 0.5 1.65
+ 26 0.5 1.675
+ 26 0.5 1.7
+ 26 0.5 1.725
+ 26 0.5 1.75
+ 26 0.5 1.775
+ 26 0.5 1.8
+ 26 0.5 1.825
+ 26 0.5 1.85
+ 26 0.5 1.875
+ 26 0.5 1.9
+ 26 0.5 1.925
+ 26 0.5 1.95
+ 26 0.5 1.975
+ 26 0.5 2.0
+ 26 0.5 2.025
+ 26 0.5 2.05
+ 26 0.5 2.075
+ 26 0.5 2.1
+ 26 0.5 2.125
+ 26 0.5 2.15
+ 26 0.5 2.175
+ 26 0.5 2.2
+ 26 0.5 2.225
+ 26 0.5 2.25
+ 26 0.5 2.275
+ 26 0.5 2.3
+ 26 0.5 2.325
+ 26 0.5 2.35
+ 26 0.5 2.375
+ 26 0.5 2.4
+ 26 0.5 2.425
+ 26 0.5 2.45
+ 26 0.5 2.475
+ 26 0.5 2.5
+ 28 0.5 1.25
+ 28 0.5 1.275
+ 28 0.5 1.3
+ 28 0.5 1.325
+ 28 0.5 1.35
+ 28 0.5 1.375
+ 28 0.5 1.4
+ 28 0.5 1.425
+ 28 0.5 1.45
+ 28 0.5 1.475
+ 28 0.5 1.5
+ 28 0.5 1.525
+ 28 0.5 1.55
+ 28 0.5 1.575
+ 28 0.5 1.6
+ 28 0.5 1.625
+ 28 0.5 1.65
+ 28 0.5 1.675
+ 28 0.5 1.7
+ 28 0.5 1.725
+ 28 0.5 1.75
+ 28 0.5 1.775
+ 28 0.5 1.8
+ 28 0.5 1.825
+ 28 0.5 1.85
+ 28 0.5 1.875
+ 28 0.5 1.9
+ 28 0.5 1.925
+ 28 0.5 1.95
+ 28 0.5 1.975
+ 28 0.5 2.0
+ 28 0.5 2.025
+ 28 0.5 2.05
+ 28 0.5 2.075
+ 28 0.5 2.1
+ 28 0.5 2.125
+ 28 0.5 2.15
+ 28 0.5 2.175
+ 28 0.5 2.2
+ 28 0.5 2.225
+ 28 0.5 2.25
+ 28 0.5 2.275
+ 28 0.5 2.3
+ 28 0.5 2.325
+ 28 0.5 2.35
+ 28 0.5 2.375
+ 28 0.5 2.4
+ 28 0.5 2.425
+ 28 0.5 2.45
+ 28 0.5 2.475
+ 28 0.5 2.5
+ 30 0.5 1.25
+ 30 0.5 1.275
+ 30 0.5 1.3
+ 30 0.5 1.325
+ 30 0.5 1.35
+ 30 0.5 1.375
+ 30 0.5 1.4
+ 30 0.5 1.425
+ 30 0.5 1.45
+ 30 0.5 1.475
+ 30 0.5 1.5
+ 30 0.5 1.525
+ 30 0.5 1.55
+ 30 0.5 1.575
+ 30 0.5 1.6
+ 30 0.5 1.625
+ 30 0.5 1.65
+ 30 0.5 1.675
+ 30 0.5 1.7
+ 30 0.5 1.725
+ 30 0.5 1.75
+ 30 0.5 1.775
+ 30 0.5 1.8
+ 30 0.5 1.825
+ 30 0.5 1.85
+ 30 0.5 1.875
+ 30 0.5 1.9
+ 30 0.5 1.925
+ 30 0.5 1.95
+ 30 0.5 1.975
+ 30 0.5 2.0
+ 30 0.5 2.025
+ 30 0.5 2.05
+ 30 0.5 2.075
+ 30 0.5 2.1
+ 30 0.5 2.125
+ 30 0.5 2.15
+ 30 0.5 2.175
+ 30 0.5 2.2
+ 30 0.5 2.225
+ 30 0.5 2.25
+ 30 0.5 2.275
+ 30 0.5 2.3
+ 30 0.5 2.325
+ 30 0.5 2.35
+ 30 0.5 2.375
+ 30 0.5 2.4
+ 30 0.5 2.425
+ 30 0.5 2.45
+ 30 0.5 2.475
+ 30 0.5 2.5
+ 32 0.5 1.25
+ 32 0.5 1.275
+ 32 0.5 1.3
+ 32 0.5 1.325
+ 32 0.5 1.35
+ 32 0.5 1.375
+ 32 0.5 1.4
+ 32 0.5 1.425
+ 32 0.5 1.45
+ 32 0.5 1.475
+ 32 0.5 1.5
+ 32 0.5 1.525
+ 32 0.5 1.55
+ 32 0.5 1.575
+ 32 0.5 1.6
+ 32 0.5 1.625
+ 32 0.5 1.65
+ 32 0.5 1.675
+ 32 0.5 1.7
+ 32 0.5 1.725
+ 32 0.5 1.75
+ 32 0.5 1.775
+ 32 0.5 1.8
+ 32 0.5 1.825
+ 32 0.5 1.85
+ 32 0.5 1.875
+ 32 0.5 1.9
+ 32 0.5 1.925
+ 32 0.5 1.95
+ 32 0.5 1.975
+ 32 0.5 2.0
+ 32 0.5 2.025
+ 32 0.5 2.05
+ 32 0.5 2.075
+ 32 0.5 2.1
+ 32 0.5 2.125
+ 32 0.5 2.15
+ 32 0.5 2.175
+ 32 0.5 2.2
+ 32 0.5 2.225
+ 32 0.5 2.25
+ 32 0.5 2.275
+ 32 0.5 2.3
+ 32 0.5 2.325
+ 32 0.5 2.35
+ 32 0.5 2.375
+ 32 0.5 2.4
+ 32 0.5 2.425
+ 32 0.5 2.45
+ 32 0.5 2.475
+ 32 0.5 2.5
+ 34 0.5 1.25
+ 34 0.5 1.275
+ 34 0.5 1.3
+ 34 0.5 1.325
+ 34 0.5 1.35
+ 34 0.5 1.375
+ 34 0.5 1.4
+ 34 0.5 1.425
+ 34 0.5 1.45
+ 34 0.5 1.475
+ 34 0.5 1.5
+ 34 0.5 1.525
+ 34 0.5 1.55
+ 34 0.5 1.575
+ 34 0.5 1.6
+ 34 0.5 1.625
+ 34 0.5 1.65
+ 34 0.5 1.675
+ 34 0.5 1.7
+ 34 0.5 1.725
+ 34 0.5 1.75
+ 34 0.5 1.775
+ 34 0.5 1.8
+ 34 0.5 1.825
+ 34 0.5 1.85
+ 34 0.5 1.875
+ 34 0.5 1.9
+ 34 0.5 1.925
+ 34 0.5 1.95
+ 34 0.5 1.975
+ 34 0.5 2.0
+ 34 0.5 2.025
+ 34 0.5 2.05
+ 34 0.5 2.075
+ 34 0.5 2.1
+ 34 0.5 2.125
+ 34 0.5 2.15
+ 34 0.5 2.175
+ 34 0.5 2.2
+ 34 0.5 2.225
+ 34 0.5 2.25
+ 34 0.5 2.275
+ 34 0.5 2.3
+ 34 0.5 2.325
+ 34 0.5 2.35
+ 34 0.5 2.375
+ 34 0.5 2.4
+ 34 0.5 2.425
+ 34 0.5 2.45
+ 34 0.5 2.475
+ 34 0.5 2.5
+ 36 0.5 1.25
+ 36 0.5 1.275
+ 36 0.5 1.3
+ 36 0.5 1.325
+ 36 0.5 1.35
+ 36 0.5 1.375
+ 36 0.5 1.4
+ 36 0.5 1.425
+ 36 0.5 1.45
+ 36 0.5 1.475
+ 36 0.5 1.5
+ 36 0.5 1.525
+ 36 0.5 1.55
+ 36 0.5 1.575
+ 36 0.5 1.6
+ 36 0.5 1.625
+ 36 0.5 1.65
+ 36 0.5 1.675
+ 36 0.5 1.7
+ 36 0.5 1.725
+ 36 0.5 1.75
+ 36 0.5 1.775
+ 36 0.5 1.8
+ 36 0.5 1.825
+ 36 0.5 1.85
+ 36 0.5 1.875
+ 36 0.5 1.9
+ 36 0.5 1.925
+ 36 0.5 1.95
+ 36 0.5 1.975
+ 36 0.5 2.0
+ 36 0.5 2.025
+ 36 0.5 2.05
+ 36 0.5 2.075
+ 36 0.5 2.1
+ 36 0.5 2.125
+ 36 0.5 2.15
+ 36 0.5 2.175
+ 36 0.5 2.2
+ 36 0.5 2.225
+ 36 0.5 2.25
+ 36 0.5 2.275
+ 36 0.5 2.3
+ 36 0.5 2.325
+ 36 0.5 2.35
+ 36 0.5 2.375
+ 36 0.5 2.4
+ 36 0.5 2.425
+ 36 0.5 2.45
+ 36 0.5 2.475
+ 36 0.5 2.5
+ 38 0.5 1.25
+ 38 0.5 1.275
+ 38 0.5 1.3
+ 38 0.5 1.325
+ 38 0.5 1.35
+ 38 0.5 1.375
+ 38 0.5 1.4
+ 38 0.5 1.425
+ 38 0.5 1.45
+ 38 0.5 1.475
+ 38 0.5 1.5
+ 38 0.5 1.525
+ 38 0.5 1.55
+ 38 0.5 1.575
+ 38 0.5 1.6
+ 38 0.5 1.625
+ 38 0.5 1.65
+ 38 0.5 1.675
+ 38 0.5 1.7
+ 38 0.5 1.725
+ 38 0.5 1.75
+ 38 0.5 1.775
+ 38 0.5 1.8
+ 38 0.5 1.825
+ 38 0.5 1.85
+ 38 0.5 1.875
+ 38 0.5 1.9
+ 38 0.5 1.925
+ 38 0.5 1.95
+ 38 0.5 1.975
+ 38 0.5 2.0
+ 38 0.5 2.025
+ 38 0.5 2.05
+ 38 0.5 2.075
+ 38 0.5 2.1
+ 38 0.5 2.125
+ 38 0.5 2.15
+ 38 0.5 2.175
+ 38 0.5 2.2
+ 38 0.5 2.225
+ 38 0.5 2.25
+ 38 0.5 2.275
+ 38 0.5 2.3
+ 38 0.5 2.325
+ 38 0.5 2.35
+ 38 0.5 2.375
+ 38 0.5 2.4
+ 38 0.5 2.425
+ 38 0.5 2.45
+ 38 0.5 2.475
+ 38 0.5 2.5
+ 40 0.5 1.25
+ 40 0.5 1.275
+ 40 0.5 1.3
+ 40 0.5 1.325
+ 40 0.5 1.35
+ 40 0.5 1.375
+ 40 0.5 1.4
+ 40 0.5 1.425
+ 40 0.5 1.45
+ 40 0.5 1.475
+ 40 0.5 1.5
+ 40 0.5 1.525
+ 40 0.5 1.55
+ 40 0.5 1.575
+ 40 0.5 1.6
+ 40 0.5 1.625
+ 40 0.5 1.65
+ 40 0.5 1.675
+ 40 0.5 1.7
+ 40 0.5 1.725
+ 40 0.5 1.75
+ 40 0.5 1.775
+ 40 0.5 1.8
+ 40 0.5 1.825
+ 40 0.5 1.85
+ 40 0.5 1.875
+ 40 0.5 1.9
+ 40 0.5 1.925
+ 40 0.5 1.95
+ 40 0.5 1.975
+ 40 0.5 2.0
+ 40 0.5 2.025
+ 40 0.5 2.05
+ 40 0.5 2.075
+ 40 0.5 2.1
+ 40 0.5 2.125
+ 40 0.5 2.15
+ 40 0.5 2.175
+ 40 0.5 2.2
+ 40 0.5 2.225
+ 40 0.5 2.25
+ 40 0.5 2.275
+ 40 0.5 2.3
+ 40 0.5 2.325
+ 40 0.5 2.35
+ 40 0.5 2.375
+ 40 0.5 2.4
+ 40 0.5 2.425
+ 40 0.5 2.45
+ 40 0.5 2.475
+ 40 0.5 2.5
+ 42 0.5 1.25
+ 42 0.5 1.275
+ 42 0.5 1.3
+ 42 0.5 1.325
+ 42 0.5 1.35
+ 42 0.5 1.375
+ 42 0.5 1.4
+ 42 0.5 1.425
+ 42 0.5 1.45
+ 42 0.5 1.475
+ 42 0.5 1.5
+ 42 0.5 1.525
+ 42 0.5 1.55
+ 42 0.5 1.575
+ 42 0.5 1.6
+ 42 0.5 1.625
+ 42 0.5 1.65
+ 42 0.5 1.675
+ 42 0.5 1.7
+ 42 0.5 1.725
+ 42 0.5 1.75
+ 42 0.5 1.775
+ 42 0.5 1.8
+ 42 0.5 1.825
+ 42 0.5 1.85
+ 42 0.5 1.875
+ 42 0.5 1.9
+ 42 0.5 1.925
+ 42 0.5 1.95
+ 42 0.5 1.975
+ 42 0.5 2.0
+ 42 0.5 2.025
+ 42 0.5 2.05
+ 42 0.5 2.075
+ 42 0.5 2.1
+ 42 0.5 2.125
+ 42 0.5 2.15
+ 42 0.5 2.175
+ 42 0.5 2.2
+ 42 0.5 2.225
+ 42 0.5 2.25
+ 42 0.5 2.275
+ 42 0.5 2.3
+ 42 0.5 2.325
+ 42 0.5 2.35
+ 42 0.5 2.375
+ 42 0.5 2.4
+ 42 0.5 2.425
+ 42 0.5 2.45
+ 42 0.5 2.475
+ 42 0.5 2.5
+ 44 0.5 1.25
+ 44 0.5 1.275
+ 44 0.5 1.3
+ 44 0.5 1.325
+ 44 0.5 1.35
+ 44 0.5 1.375
+ 44 0.5 1.4
+ 44 0.5 1.425
+ 44 0.5 1.45
+ 44 0.5 1.475
+ 44 0.5 1.5
+ 44 0.5 1.525
+ 44 0.5 1.55
+ 44 0.5 1.575
+ 44 0.5 1.6
+ 44 0.5 1.625
+ 44 0.5 1.65
+ 44 0.5 1.675
+ 44 0.5 1.7
+ 44 0.5 1.725
+ 44 0.5 1.75
+ 44 0.5 1.775
+ 44 0.5 1.8
+ 44 0.5 1.825
+ 44 0.5 1.85
+ 44 0.5 1.875
+ 44 0.5 1.9
+ 44 0.5 1.925
+ 44 0.5 1.95
+ 44 0.5 1.975
+ 44 0.5 2.0
+ 44 0.5 2.025
+ 44 0.5 2.05
+ 44 0.5 2.075
+ 44 0.5 2.1
+ 44 0.5 2.125
+ 44 0.5 2.15
+ 44 0.5 2.175
+ 44 0.5 2.2
+ 44 0.5 2.225
+ 44 0.5 2.25
+ 44 0.5 2.275
+ 44 0.5 2.3
+ 44 0.5 2.325
+ 44 0.5 2.35
+ 44 0.5 2.375
+ 44 0.5 2.4
+ 44 0.5 2.425
+ 44 0.5 2.45
+ 44 0.5 2.475
+ 44 0.5 2.5
+ 46 0.5 1.25
+ 46 0.5 1.275
+ 46 0.5 1.3
+ 46 0.5 1.325
+ 46 0.5 1.35
+ 46 0.5 1.375
+ 46 0.5 1.4
+ 46 0.5 1.425
+ 46 0.5 1.45
+ 46 0.5 1.475
+ 46 0.5 1.5
+ 46 0.5 1.525
+ 46 0.5 1.55
+ 46 0.5 1.575
+ 46 0.5 1.6
+ 46 0.5 1.625
+ 46 0.5 1.65
+ 46 0.5 1.675
+ 46 0.5 1.7
+ 46 0.5 1.725
+ 46 0.5 1.75
+ 46 0.5 1.775
+ 46 0.5 1.8
+ 46 0.5 1.825
+ 46 0.5 1.85
+ 46 0.5 1.875
+ 46 0.5 1.9
+ 46 0.5 1.925
+ 46 0.5 1.95
+ 46 0.5 1.975
+ 46 0.5 2.0
+ 46 0.5 2.025
+ 46 0.5 2.05
+ 46 0.5 2.075
+ 46 0.5 2.1
+ 46 0.5 2.125
+ 46 0.5 2.15
+ 46 0.5 2.175
+ 46 0.5 2.2
+ 46 0.5 2.225
+ 46 0.5 2.25
+ 46 0.5 2.275
+ 46 0.5 2.3
+ 46 0.5 2.325
+ 46 0.5 2.35
+ 46 0.5 2.375
+ 46 0.5 2.4
+ 46 0.5 2.425
+ 46 0.5 2.45
+ 46 0.5 2.475
+ 46 0.5 2.5
+ 48 0.5 1.25
+ 48 0.5 1.275
+ 48 0.5 1.3
+ 48 0.5 1.325
+ 48 0.5 1.35
+ 48 0.5 1.375
+ 48 0.5 1.4
+ 48 0.5 1.425
+ 48 0.5 1.45
+ 48 0.5 1.475
+ 48 0.5 1.5
+ 48 0.5 1.525
+ 48 0.5 1.55
+ 48 0.5 1.575
+ 48 0.5 1.6
+ 48 0.5 1.625
+ 48 0.5 1.65
+ 48 0.5 1.675
+ 48 0.5 1.7
+ 48 0.5 1.725
+ 48 0.5 1.75
+ 48 0.5 1.775
+ 48 0.5 1.8
+ 48 0.5 1.825
+ 48 0.5 1.85
+ 48 0.5 1.875
+ 48 0.5 1.9
+ 48 0.5 1.925
+ 48 0.5 1.95
+ 48 0.5 1.975
+ 48 0.5 2.0
+ 48 0.5 2.025
+ 48 0.5 2.05
+ 48 0.5 2.075
+ 48 0.5 2.1
+ 48 0.5 2.125
+ 48 0.5 2.15
+ 48 0.5 2.175
+ 48 0.5 2.2
+ 48 0.5 2.225
+ 48 0.5 2.25
+ 48 0.5 2.275
+ 48 0.5 2.3
+ 48 0.5 2.325
+ 48 0.5 2.35
+ 48 0.5 2.375
+ 48 0.5 2.4
+ 48 0.5 2.425
+ 48 0.5 2.45
+ 48 0.5 2.475
+ 48 0.5 2.5
+ 50 0.5 1.25
+ 50 0.5 1.275
+ 50 0.5 1.3
+ 50 0.5 1.325
+ 50 0.5 1.35
+ 50 0.5 1.375
+ 50 0.5 1.4
+ 50 0.5 1.425
+ 50 0.5 1.45
+ 50 0.5 1.475
+ 50 0.5 1.5
+ 50 0.5 1.525
+ 50 0.5 1.55
+ 50 0.5 1.575
+ 50 0.5 1.6
+ 50 0.5 1.625
+ 50 0.5 1.65
+ 50 0.5 1.675
+ 50 0.5 1.7
+ 50 0.5 1.725
+ 50 0.5 1.75
+ 50 0.5 1.775
+ 50 0.5 1.8
+ 50 0.5 1.825
+ 50 0.5 1.85
+ 50 0.5 1.875
+ 50 0.5 1.9
+ 50 0.5 1.925
+ 50 0.5 1.95
+ 50 0.5 1.975
+ 50 0.5 2.0
+ 50 0.5 2.025
+ 50 0.5 2.05
+ 50 0.5 2.075
+ 50 0.5 2.1
+ 50 0.5 2.125
+ 50 0.5 2.15
+ 50 0.5 2.175
+ 50 0.5 2.2
+ 50 0.5 2.225
+ 50 0.5 2.25
+ 50 0.5 2.275
+ 50 0.5 2.3
+ 50 0.5 2.325
+ 50 0.5 2.35
+ 50 0.5 2.375
+ 50 0.5 2.4
+ 50 0.5 2.425
+ 50 0.5 2.45
+ 50 0.5 2.475
+ 50 0.5 2.5
+ 52 0.5 1.25
+ 52 0.5 1.275
+ 52 0.5 1.3
+ 52 0.5 1.325
+ 52 0.5 1.35
+ 52 0.5 1.375
+ 52 0.5 1.4
+ 52 0.5 1.425
+ 52 0.5 1.45
+ 52 0.5 1.475
+ 52 0.5 1.5
+ 52 0.5 1.525
+ 52 0.5 1.55
+ 52 0.5 1.575
+ 52 0.5 1.6
+ 52 0.5 1.625
+ 52 0.5 1.65
+ 52 0.5 1.675
+ 52 0.5 1.7
+ 52 0.5 1.725
+ 52 0.5 1.75
+ 52 0.5 1.775
+ 52 0.5 1.8
+ 52 0.5 1.825
+ 52 0.5 1.85
+ 52 0.5 1.875
+ 52 0.5 1.9
+ 52 0.5 1.925
+ 52 0.5 1.95
+ 52 0.5 1.975
+ 52 0.5 2.0
+ 52 0.5 2.025
+ 52 0.5 2.05
+ 52 0.5 2.075
+ 52 0.5 2.1
+ 52 0.5 2.125
+ 52 0.5 2.15
+ 52 0.5 2.175
+ 52 0.5 2.2
+ 52 0.5 2.225
+ 52 0.5 2.25
+ 52 0.5 2.275
+ 52 0.5 2.3
+ 52 0.5 2.325
+ 52 0.5 2.35
+ 52 0.5 2.375
+ 52 0.5 2.4
+ 52 0.5 2.425
+ 52 0.5 2.45
+ 52 0.5 2.475
+ 52 0.5 2.5
+ 54 0.5 1.25
+ 54 0.5 1.275
+ 54 0.5 1.3
+ 54 0.5 1.325
+ 54 0.5 1.35
+ 54 0.5 1.375
+ 54 0.5 1.4
+ 54 0.5 1.425
+ 54 0.5 1.45
+ 54 0.5 1.475
+ 54 0.5 1.5
+ 54 0.5 1.525
+ 54 0.5 1.55
+ 54 0.5 1.575
+ 54 0.5 1.6
+ 54 0.5 1.625
+ 54 0.5 1.65
+ 54 0.5 1.675
+ 54 0.5 1.7
+ 54 0.5 1.725
+ 54 0.5 1.75
+ 54 0.5 1.775
+ 54 0.5 1.8
+ 54 0.5 1.825
+ 54 0.5 1.85
+ 54 0.5 1.875
+ 54 0.5 1.9
+ 54 0.5 1.925
+ 54 0.5 1.95
+ 54 0.5 1.975
+ 54 0.5 2.0
+ 54 0.5 2.025
+ 54 0.5 2.05
+ 54 0.5 2.075
+ 54 0.5 2.1
+ 54 0.5 2.125
+ 54 0.5 2.15
+ 54 0.5 2.175
+ 54 0.5 2.2
+ 54 0.5 2.225
+ 54 0.5 2.25
+ 54 0.5 2.275
+ 54 0.5 2.3
+ 54 0.5 2.325
+ 54 0.5 2.35
+ 54 0.5 2.375
+ 54 0.5 2.4
+ 54 0.5 2.425
+ 54 0.5 2.45
+ 54 0.5 2.475
+ 54 0.5 2.5
+ 56 0.5 1.25
+ 56 0.5 1.275
+ 56 0.5 1.3
+ 56 0.5 1.325
+ 56 0.5 1.35
+ 56 0.5 1.375
+ 56 0.5 1.4
+ 56 0.5 1.425
+ 56 0.5 1.45
+ 56 0.5 1.475
+ 56 0.5 1.5
+ 56 0.5 1.525
+ 56 0.5 1.55
+ 56 0.5 1.575
+ 56 0.5 1.6
+ 56 0.5 1.625
+ 56 0.5 1.65
+ 56 0.5 1.675
+ 56 0.5 1.7
+ 56 0.5 1.725
+ 56 0.5 1.75
+ 56 0.5 1.775
+ 56 0.5 1.8
+ 56 0.5 1.825
+ 56 0.5 1.85
+ 56 0.5 1.875
+ 56 0.5 1.9
+ 56 0.5 1.925
+ 56 0.5 1.95
+ 56 0.5 1.975
+ 56 0.5 2.0
+ 56 0.5 2.025
+ 56 0.5 2.05
+ 56 0.5 2.075
+ 56 0.5 2.1
+ 56 0.5 2.125
+ 56 0.5 2.15
+ 56 0.5 2.175
+ 56 0.5 2.2
+ 56 0.5 2.225
+ 56 0.5 2.25
+ 56 0.5 2.275
+ 56 0.5 2.3
+ 56 0.5 2.325
+ 56 0.5 2.35
+ 56 0.5 2.375
+ 56 0.5 2.4
+ 56 0.5 2.425
+ 56 0.5 2.45
+ 56 0.5 2.475
+ 56 0.5 2.5
+ 58 0.5 1.25
+ 58 0.5 1.275
+ 58 0.5 1.3
+ 58 0.5 1.325
+ 58 0.5 1.35
+ 58 0.5 1.375
+ 58 0.5 1.4
+ 58 0.5 1.425
+ 58 0.5 1.45
+ 58 0.5 1.475
+ 58 0.5 1.5
+ 58 0.5 1.525
+ 58 0.5 1.55
+ 58 0.5 1.575
+ 58 0.5 1.6
+ 58 0.5 1.625
+ 58 0.5 1.65
+ 58 0.5 1.675
+ 58 0.5 1.7
+ 58 0.5 1.725
+ 58 0.5 1.75
+ 58 0.5 1.775
+ 58 0.5 1.8
+ 58 0.5 1.825
+ 58 0.5 1.85
+ 58 0.5 1.875
+ 58 0.5 1.9
+ 58 0.5 1.925
+ 58 0.5 1.95
+ 58 0.5 1.975
+ 58 0.5 2.0
+ 58 0.5 2.025
+ 58 0.5 2.05
+ 58 0.5 2.075
+ 58 0.5 2.1
+ 58 0.5 2.125
+ 58 0.5 2.15
+ 58 0.5 2.175
+ 58 0.5 2.2
+ 58 0.5 2.225
+ 58 0.5 2.25
+ 58 0.5 2.275
+ 58 0.5 2.3
+ 58 0.5 2.325
+ 58 0.5 2.35
+ 58 0.5 2.375
+ 58 0.5 2.4
+ 58 0.5 2.425
+ 58 0.5 2.45
+ 58 0.5 2.475
+ 58 0.5 2.5
+ 60 0.5 1.25
+ 60 0.5 1.275
+ 60 0.5 1.3
+ 60 0.5 1.325
+ 60 0.5 1.35
+ 60 0.5 1.375
+ 60 0.5 1.4
+ 60 0.5 1.425
+ 60 0.5 1.45
+ 60 0.5 1.475
+ 60 0.5 1.5
+ 60 0.5 1.525
+ 60 0.5 1.55
+ 60 0.5 1.575
+ 60 0.5 1.6
+ 60 0.5 1.625
+ 60 0.5 1.65
+ 60 0.5 1.675
+ 60 0.5 1.7
+ 60 0.5 1.725
+ 60 0.5 1.75
+ 60 0.5 1.775
+ 60 0.5 1.8
+ 60 0.5 1.825
+ 60 0.5 1.85
+ 60 0.5 1.875
+ 60 0.5 1.9
+ 60 0.5 1.925
+ 60 0.5 1.95
+ 60 0.5 1.975
+ 60 0.5 2.0
+ 60 0.5 2.025
+ 60 0.5 2.05
+ 60 0.5 2.075
+ 60 0.5 2.1
+ 60 0.5 2.125
+ 60 0.5 2.15
+ 60 0.5 2.175
+ 60 0.5 2.2
+ 60 0.5 2.225
+ 60 0.5 2.25
+ 60 0.5 2.275
+ 60 0.5 2.3
+ 60 0.5 2.325
+ 60 0.5 2.35
+ 60 0.5 2.375
+ 60 0.5 2.4
+ 60 0.5 2.425
+ 60 0.5 2.45
+ 60 0.5 2.475
+ 60 0.5 2.5
+ 62 0.5 1.25
+ 62 0.5 1.275
+ 62 0.5 1.3
+ 62 0.5 1.325
+ 62 0.5 1.35
+ 62 0.5 1.375
+ 62 0.5 1.4
+ 62 0.5 1.425
+ 62 0.5 1.45
+ 62 0.5 1.475
+ 62 0.5 1.5
+ 62 0.5 1.525
+ 62 0.5 1.55
+ 62 0.5 1.575
+ 62 0.5 1.6
+ 62 0.5 1.625
+ 62 0.5 1.65
+ 62 0.5 1.675
+ 62 0.5 1.7
+ 62 0.5 1.725
+ 62 0.5 1.75
+ 62 0.5 1.775
+ 62 0.5 1.8
+ 62 0.5 1.825
+ 62 0.5 1.85
+ 62 0.5 1.875
+ 62 0.5 1.9
+ 62 0.5 1.925
+ 62 0.5 1.95
+ 62 0.5 1.975
+ 62 0.5 2.0
+ 62 0.5 2.025
+ 62 0.5 2.05
+ 62 0.5 2.075
+ 62 0.5 2.1
+ 62 0.5 2.125
+ 62 0.5 2.15
+ 62 0.5 2.175
+ 62 0.5 2.2
+ 62 0.5 2.225
+ 62 0.5 2.25
+ 62 0.5 2.275
+ 62 0.5 2.3
+ 62 0.5 2.325
+ 62 0.5 2.35
+ 62 0.5 2.375
+ 62 0.5 2.4
+ 62 0.5 2.425
+ 62 0.5 2.45
+ 62 0.5 2.475
+ 62 0.5 2.5
+ 64 0.5 1.25
+ 64 0.5 1.275
+ 64 0.5 1.3
+ 64 0.5 1.325
+ 64 0.5 1.35
+ 64 0.5 1.375
+ 64 0.5 1.4
+ 64 0.5 1.425
+ 64 0.5 1.45
+ 64 0.5 1.475
+ 64 0.5 1.5
+ 64 0.5 1.525
+ 64 0.5 1.55
+ 64 0.5 1.575
+ 64 0.5 1.6
+ 64 0.5 1.625
+ 64 0.5 1.65
+ 64 0.5 1.675
+ 64 0.5 1.7
+ 64 0.5 1.725
+ 64 0.5 1.75
+ 64 0.5 1.775
+ 64 0.5 1.8
+ 64 0.5 1.825
+ 64 0.5 1.85
+ 64 0.5 1.875
+ 64 0.5 1.9
+ 64 0.5 1.925
+ 64 0.5 1.95
+ 64 0.5 1.975
+ 64 0.5 2.0
+ 64 0.5 2.025
+ 64 0.5 2.05
+ 64 0.5 2.075
+ 64 0.5 2.1
+ 64 0.5 2.125
+ 64 0.5 2.15
+ 64 0.5 2.175
+ 64 0.5 2.2
+ 64 0.5 2.225
+ 64 0.5 2.25
+ 64 0.5 2.275
+ 64 0.5 2.3
+ 64 0.5 2.325
+ 64 0.5 2.35
+ 64 0.5 2.375
+ 64 0.5 2.4
+ 64 0.5 2.425
+ 64 0.5 2.45
+ 64 0.5 2.475
+ 64 0.5 2.5
+ 66 0.5 1.25
+ 66 0.5 1.275
+ 66 0.5 1.3
+ 66 0.5 1.325
+ 66 0.5 1.35
+ 66 0.5 1.375
+ 66 0.5 1.4
+ 66 0.5 1.425
+ 66 0.5 1.45
+ 66 0.5 1.475
+ 66 0.5 1.5
+ 66 0.5 1.525
+ 66 0.5 1.55
+ 66 0.5 1.575
+ 66 0.5 1.6
+ 66 0.5 1.625
+ 66 0.5 1.65
+ 66 0.5 1.675
+ 66 0.5 1.7
+ 66 0.5 1.725
+ 66 0.5 1.75
+ 66 0.5 1.775
+ 66 0.5 1.8
+ 66 0.5 1.825
+ 66 0.5 1.85
+ 66 0.5 1.875
+ 66 0.5 1.9
+ 66 0.5 1.925
+ 66 0.5 1.95
+ 66 0.5 1.975
+ 66 0.5 2.0
+ 66 0.5 2.025
+ 66 0.5 2.05
+ 66 0.5 2.075
+ 66 0.5 2.1
+ 66 0.5 2.125
+ 66 0.5 2.15
+ 66 0.5 2.175
+ 66 0.5 2.2
+ 66 0.5 2.225
+ 66 0.5 2.25
+ 66 0.5 2.275
+ 66 0.5 2.3
+ 66 0.5 2.325
+ 66 0.5 2.35
+ 66 0.5 2.375
+ 66 0.5 2.4
+ 66 0.5 2.425
+ 66 0.5 2.45
+ 66 0.5 2.475
+ 66 0.5 2.5
+ 68 0.5 1.25
+ 68 0.5 1.275
+ 68 0.5 1.3
+ 68 0.5 1.325
+ 68 0.5 1.35
+ 68 0.5 1.375
+ 68 0.5 1.4
+ 68 0.5 1.425
+ 68 0.5 1.45
+ 68 0.5 1.475
+ 68 0.5 1.5
+ 68 0.5 1.525
+ 68 0.5 1.55
+ 68 0.5 1.575
+ 68 0.5 1.6
+ 68 0.5 1.625
+ 68 0.5 1.65
+ 68 0.5 1.675
+ 68 0.5 1.7
+ 68 0.5 1.725
+ 68 0.5 1.75
+ 68 0.5 1.775
+ 68 0.5 1.8
+ 68 0.5 1.825
+ 68 0.5 1.85
+ 68 0.5 1.875
+ 68 0.5 1.9
+ 68 0.5 1.925
+ 68 0.5 1.95
+ 68 0.5 1.975
+ 68 0.5 2.0
+ 68 0.5 2.025
+ 68 0.5 2.05
+ 68 0.5 2.075
+ 68 0.5 2.1
+ 68 0.5 2.125
+ 68 0.5 2.15
+ 68 0.5 2.175
+ 68 0.5 2.2
+ 68 0.5 2.225
+ 68 0.5 2.25
+ 68 0.5 2.275
+ 68 0.5 2.3
+ 68 0.5 2.325
+ 68 0.5 2.35
+ 68 0.5 2.375
+ 68 0.5 2.4
+ 68 0.5 2.425
+ 68 0.5 2.45
+ 68 0.5 2.475
+ 68 0.5 2.5
+ 70 0.5 1.25
+ 70 0.5 1.275
+ 70 0.5 1.3
+ 70 0.5 1.325
+ 70 0.5 1.35
+ 70 0.5 1.375
+ 70 0.5 1.4
+ 70 0.5 1.425
+ 70 0.5 1.45
+ 70 0.5 1.475
+ 70 0.5 1.5
+ 70 0.5 1.525
+ 70 0.5 1.55
+ 70 0.5 1.575
+ 70 0.5 1.6
+ 70 0.5 1.625
+ 70 0.5 1.65
+ 70 0.5 1.675
+ 70 0.5 1.7
+ 70 0.5 1.725
+ 70 0.5 1.75
+ 70 0.5 1.775
+ 70 0.5 1.8
+ 70 0.5 1.825
+ 70 0.5 1.85
+ 70 0.5 1.875
+ 70 0.5 1.9
+ 70 0.5 1.925
+ 70 0.5 1.95
+ 70 0.5 1.975
+ 70 0.5 2.0
+ 70 0.5 2.025
+ 70 0.5 2.05
+ 70 0.5 2.075
+ 70 0.5 2.1
+ 70 0.5 2.125
+ 70 0.5 2.15
+ 70 0.5 2.175
+ 70 0.5 2.2
+ 70 0.5 2.225
+ 70 0.5 2.25
+ 70 0.5 2.275
+ 70 0.5 2.3
+ 70 0.5 2.325
+ 70 0.5 2.35
+ 70 0.5 2.375
+ 70 0.5 2.4
+ 70 0.5 2.425
+ 70 0.5 2.45
+ 70 0.5 2.475
+ 70 0.5 2.5
+ 72 0.5 1.25
+ 72 0.5 1.275
+ 72 0.5 1.3
+ 72 0.5 1.325
+ 72 0.5 1.35
+ 72 0.5 1.375
+ 72 0.5 1.4
+ 72 0.5 1.425
+ 72 0.5 1.45
+ 72 0.5 1.475
+ 72 0.5 1.5
+ 72 0.5 1.525
+ 72 0.5 1.55
+ 72 0.5 1.575
+ 72 0.5 1.6
+ 72 0.5 1.625
+ 72 0.5 1.65
+ 72 0.5 1.675
+ 72 0.5 1.7
+ 72 0.5 1.725
+ 72 0.5 1.75
+ 72 0.5 1.775
+ 72 0.5 1.8
+ 72 0.5 1.825
+ 72 0.5 1.85
+ 72 0.5 1.875
+ 72 0.5 1.9
+ 72 0.5 1.925
+ 72 0.5 1.95
+ 72 0.5 1.975
+ 72 0.5 2.0
+ 72 0.5 2.025
+ 72 0.5 2.05
+ 72 0.5 2.075
+ 72 0.5 2.1
+ 72 0.5 2.125
+ 72 0.5 2.15
+ 72 0.5 2.175
+ 72 0.5 2.2
+ 72 0.5 2.225
+ 72 0.5 2.25
+ 72 0.5 2.275
+ 72 0.5 2.3
+ 72 0.5 2.325
+ 72 0.5 2.35
+ 72 0.5 2.375
+ 72 0.5 2.4
+ 72 0.5 2.425
+ 72 0.5 2.45
+ 72 0.5 2.475
+ 72 0.5 2.5
+ 74 0.5 1.25
+ 74 0.5 1.275
+ 74 0.5 1.3
+ 74 0.5 1.325
+ 74 0.5 1.35
+ 74 0.5 1.375
+ 74 0.5 1.4
+ 74 0.5 1.425
+ 74 0.5 1.45
+ 74 0.5 1.475
+ 74 0.5 1.5
+ 74 0.5 1.525
+ 74 0.5 1.55
+ 74 0.5 1.575
+ 74 0.5 1.6
+ 74 0.5 1.625
+ 74 0.5 1.65
+ 74 0.5 1.675
+ 74 0.5 1.7
+ 74 0.5 1.725
+ 74 0.5 1.75
+ 74 0.5 1.775
+ 74 0.5 1.8
+ 74 0.5 1.825
+ 74 0.5 1.85
+ 74 0.5 1.875
+ 74 0.5 1.9
+ 74 0.5 1.925
+ 74 0.5 1.95
+ 74 0.5 1.975
+ 74 0.5 2.0
+ 74 0.5 2.025
+ 74 0.5 2.05
+ 74 0.5 2.075
+ 74 0.5 2.1
+ 74 0.5 2.125
+ 74 0.5 2.15
+ 74 0.5 2.175
+ 74 0.5 2.2
+ 74 0.5 2.225
+ 74 0.5 2.25
+ 74 0.5 2.275
+ 74 0.5 2.3
+ 74 0.5 2.325
+ 74 0.5 2.35
+ 74 0.5 2.375
+ 74 0.5 2.4
+ 74 0.5 2.425
+ 74 0.5 2.45
+ 74 0.5 2.475
+ 74 0.5 2.5
+ 76 0.5 1.25
+ 76 0.5 1.275
+ 76 0.5 1.3
+ 76 0.5 1.325
+ 76 0.5 1.35
+ 76 0.5 1.375
+ 76 0.5 1.4
+ 76 0.5 1.425
+ 76 0.5 1.45
+ 76 0.5 1.475
+ 76 0.5 1.5
+ 76 0.5 1.525
+ 76 0.5 1.55
+ 76 0.5 1.575
+ 76 0.5 1.6
+ 76 0.5 1.625
+ 76 0.5 1.65
+ 76 0.5 1.675
+ 76 0.5 1.7
+ 76 0.5 1.725
+ 76 0.5 1.75
+ 76 0.5 1.775
+ 76 0.5 1.8
+ 76 0.5 1.825
+ 76 0.5 1.85
+ 76 0.5 1.875
+ 76 0.5 1.9
+ 76 0.5 1.925
+ 76 0.5 1.95
+ 76 0.5 1.975
+ 76 0.5 2.0
+ 76 0.5 2.025
+ 76 0.5 2.05
+ 76 0.5 2.075
+ 76 0.5 2.1
+ 76 0.5 2.125
+ 76 0.5 2.15
+ 76 0.5 2.175
+ 76 0.5 2.2
+ 76 0.5 2.225
+ 76 0.5 2.25
+ 76 0.5 2.275
+ 76 0.5 2.3
+ 76 0.5 2.325
+ 76 0.5 2.35
+ 76 0.5 2.375
+ 76 0.5 2.4
+ 76 0.5 2.425
+ 76 0.5 2.45
+ 76 0.5 2.475
+ 76 0.5 2.5
+ 78 0.5 1.25
+ 78 0.5 1.275
+ 78 0.5 1.3
+ 78 0.5 1.325
+ 78 0.5 1.35
+ 78 0.5 1.375
+ 78 0.5 1.4
+ 78 0.5 1.425
+ 78 0.5 1.45
+ 78 0.5 1.475
+ 78 0.5 1.5
+ 78 0.5 1.525
+ 78 0.5 1.55
+ 78 0.5 1.575
+ 78 0.5 1.6
+ 78 0.5 1.625
+ 78 0.5 1.65
+ 78 0.5 1.675
+ 78 0.5 1.7
+ 78 0.5 1.725
+ 78 0.5 1.75
+ 78 0.5 1.775
+ 78 0.5 1.8
+ 78 0.5 1.825
+ 78 0.5 1.85
+ 78 0.5 1.875
+ 78 0.5 1.9
+ 78 0.5 1.925
+ 78 0.5 1.95
+ 78 0.5 1.975
+ 78 0.5 2.0
+ 78 0.5 2.025
+ 78 0.5 2.05
+ 78 0.5 2.075
+ 78 0.5 2.1
+ 78 0.5 2.125
+ 78 0.5 2.15
+ 78 0.5 2.175
+ 78 0.5 2.2
+ 78 0.5 2.225
+ 78 0.5 2.25
+ 78 0.5 2.275
+ 78 0.5 2.3
+ 78 0.5 2.325
+ 78 0.5 2.35
+ 78 0.5 2.375
+ 78 0.5 2.4
+ 78 0.5 2.425
+ 78 0.5 2.45
+ 78 0.5 2.475
+ 78 0.5 2.5
+ 80 0.5 1.25
+ 80 0.5 1.275
+ 80 0.5 1.3
+ 80 0.5 1.325
+ 80 0.5 1.35
+ 80 0.5 1.375
+ 80 0.5 1.4
+ 80 0.5 1.425
+ 80 0.5 1.45
+ 80 0.5 1.475
+ 80 0.5 1.5
+ 80 0.5 1.525
+ 80 0.5 1.55
+ 80 0.5 1.575
+ 80 0.5 1.6
+ 80 0.5 1.625
+ 80 0.5 1.65
+ 80 0.5 1.675
+ 80 0.5 1.7
+ 80 0.5 1.725
+ 80 0.5 1.75
+ 80 0.5 1.775
+ 80 0.5 1.8
+ 80 0.5 1.825
+ 80 0.5 1.85
+ 80 0.5 1.875
+ 80 0.5 1.9
+ 80 0.5 1.925
+ 80 0.5 1.95
+ 80 0.5 1.975
+ 80 0.5 2.0
+ 80 0.5 2.025
+ 80 0.5 2.05
+ 80 0.5 2.075
+ 80 0.5 2.1
+ 80 0.5 2.125
+ 80 0.5 2.15
+ 80 0.5 2.175
+ 80 0.5 2.2
+ 80 0.5 2.225
+ 80 0.5 2.25
+ 80 0.5 2.275
+ 80 0.5 2.3
+ 80 0.5 2.325
+ 80 0.5 2.35
+ 80 0.5 2.375
+ 80 0.5 2.4
+ 80 0.5 2.425
+ 80 0.5 2.45
+ 80 0.5 2.475
+ 80 0.5 2.5
+ 82 0.5 1.25
+ 82 0.5 1.275
+ 82 0.5 1.3
+ 82 0.5 1.325
+ 82 0.5 1.35
+ 82 0.5 1.375
+ 82 0.5 1.4
+ 82 0.5 1.425
+ 82 0.5 1.45
+ 82 0.5 1.475
+ 82 0.5 1.5
+ 82 0.5 1.525
+ 82 0.5 1.55
+ 82 0.5 1.575
+ 82 0.5 1.6
+ 82 0.5 1.625
+ 82 0.5 1.65
+ 82 0.5 1.675
+ 82 0.5 1.7
+ 82 0.5 1.725
+ 82 0.5 1.75
+ 82 0.5 1.775
+ 82 0.5 1.8
+ 82 0.5 1.825
+ 82 0.5 1.85
+ 82 0.5 1.875
+ 82 0.5 1.9
+ 82 0.5 1.925
+ 82 0.5 1.95
+ 82 0.5 1.975
+ 82 0.5 2.0
+ 82 0.5 2.025
+ 82 0.5 2.05
+ 82 0.5 2.075
+ 82 0.5 2.1
+ 82 0.5 2.125
+ 82 0.5 2.15
+ 82 0.5 2.175
+ 82 0.5 2.2
+ 82 0.5 2.225
+ 82 0.5 2.25
+ 82 0.5 2.275
+ 82 0.5 2.3
+ 82 0.5 2.325
+ 82 0.5 2.35
+ 82 0.5 2.375
+ 82 0.5 2.4
+ 82 0.5 2.425
+ 82 0.5 2.45
+ 82 0.5 2.475
+ 82 0.5 2.5
+ 84 0.5 1.25
+ 84 0.5 1.275
+ 84 0.5 1.3
+ 84 0.5 1.325
+ 84 0.5 1.35
+ 84 0.5 1.375
+ 84 0.5 1.4
+ 84 0.5 1.425
+ 84 0.5 1.45
+ 84 0.5 1.475
+ 84 0.5 1.5
+ 84 0.5 1.525
+ 84 0.5 1.55
+ 84 0.5 1.575
+ 84 0.5 1.6
+ 84 0.5 1.625
+ 84 0.5 1.65
+ 84 0.5 1.675
+ 84 0.5 1.7
+ 84 0.5 1.725
+ 84 0.5 1.75
+ 84 0.5 1.775
+ 84 0.5 1.8
+ 84 0.5 1.825
+ 84 0.5 1.85
+ 84 0.5 1.875
+ 84 0.5 1.9
+ 84 0.5 1.925
+ 84 0.5 1.95
+ 84 0.5 1.975
+ 84 0.5 2.0
+ 84 0.5 2.025
+ 84 0.5 2.05
+ 84 0.5 2.075
+ 84 0.5 2.1
+ 84 0.5 2.125
+ 84 0.5 2.15
+ 84 0.5 2.175
+ 84 0.5 2.2
+ 84 0.5 2.225
+ 84 0.5 2.25
+ 84 0.5 2.275
+ 84 0.5 2.3
+ 84 0.5 2.325
+ 84 0.5 2.35
+ 84 0.5 2.375
+ 84 0.5 2.4
+ 84 0.5 2.425
+ 84 0.5 2.45
+ 84 0.5 2.475
+ 84 0.5 2.5
+ 86 0.5 1.25
+ 86 0.5 1.275
+ 86 0.5 1.3
+ 86 0.5 1.325
+ 86 0.5 1.35
+ 86 0.5 1.375
+ 86 0.5 1.4
+ 86 0.5 1.425
+ 86 0.5 1.45
+ 86 0.5 1.475
+ 86 0.5 1.5
+ 86 0.5 1.525
+ 86 0.5 1.55
+ 86 0.5 1.575
+ 86 0.5 1.6
+ 86 0.5 1.625
+ 86 0.5 1.65
+ 86 0.5 1.675
+ 86 0.5 1.7
+ 86 0.5 1.725
+ 86 0.5 1.75
+ 86 0.5 1.775
+ 86 0.5 1.8
+ 86 0.5 1.825
+ 86 0.5 1.85
+ 86 0.5 1.875
+ 86 0.5 1.9
+ 86 0.5 1.925
+ 86 0.5 1.95
+ 86 0.5 1.975
+ 86 0.5 2.0
+ 86 0.5 2.025
+ 86 0.5 2.05
+ 86 0.5 2.075
+ 86 0.5 2.1
+ 86 0.5 2.125
+ 86 0.5 2.15
+ 86 0.5 2.175
+ 86 0.5 2.2
+ 86 0.5 2.225
+ 86 0.5 2.25
+ 86 0.5 2.275
+ 86 0.5 2.3
+ 86 0.5 2.325
+ 86 0.5 2.35
+ 86 0.5 2.375
+ 86 0.5 2.4
+ 86 0.5 2.425
+ 86 0.5 2.45
+ 86 0.5 2.475
+ 86 0.5 2.5
+ 88 0.5 1.25
+ 88 0.5 1.275
+ 88 0.5 1.3
+ 88 0.5 1.325
+ 88 0.5 1.35
+ 88 0.5 1.375
+ 88 0.5 1.4
+ 88 0.5 1.425
+ 88 0.5 1.45
+ 88 0.5 1.475
+ 88 0.5 1.5
+ 88 0.5 1.525
+ 88 0.5 1.55
+ 88 0.5 1.575
+ 88 0.5 1.6
+ 88 0.5 1.625
+ 88 0.5 1.65
+ 88 0.5 1.675
+ 88 0.5 1.7
+ 88 0.5 1.725
+ 88 0.5 1.75
+ 88 0.5 1.775
+ 88 0.5 1.8
+ 88 0.5 1.825
+ 88 0.5 1.85
+ 88 0.5 1.875
+ 88 0.5 1.9
+ 88 0.5 1.925
+ 88 0.5 1.95
+ 88 0.5 1.975
+ 88 0.5 2.0
+ 88 0.5 2.025
+ 88 0.5 2.05
+ 88 0.5 2.075
+ 88 0.5 2.1
+ 88 0.5 2.125
+ 88 0.5 2.15
+ 88 0.5 2.175
+ 88 0.5 2.2
+ 88 0.5 2.225
+ 88 0.5 2.25
+ 88 0.5 2.275
+ 88 0.5 2.3
+ 88 0.5 2.325
+ 88 0.5 2.35
+ 88 0.5 2.375
+ 88 0.5 2.4
+ 88 0.5 2.425
+ 88 0.5 2.45
+ 88 0.5 2.475
+ 88 0.5 2.5
+ 90 0.5 1.25
+ 90 0.5 1.275
+ 90 0.5 1.3
+ 90 0.5 1.325
+ 90 0.5 1.35
+ 90 0.5 1.375
+ 90 0.5 1.4
+ 90 0.5 1.425
+ 90 0.5 1.45
+ 90 0.5 1.475
+ 90 0.5 1.5
+ 90 0.5 1.525
+ 90 0.5 1.55
+ 90 0.5 1.575
+ 90 0.5 1.6
+ 90 0.5 1.625
+ 90 0.5 1.65
+ 90 0.5 1.675
+ 90 0.5 1.7
+ 90 0.5 1.725
+ 90 0.5 1.75
+ 90 0.5 1.775
+ 90 0.5 1.8
+ 90 0.5 1.825
+ 90 0.5 1.85
+ 90 0.5 1.875
+ 90 0.5 1.9
+ 90 0.5 1.925
+ 90 0.5 1.95
+ 90 0.5 1.975
+ 90 0.5 2.0
+ 90 0.5 2.025
+ 90 0.5 2.05
+ 90 0.5 2.075
+ 90 0.5 2.1
+ 90 0.5 2.125
+ 90 0.5 2.15
+ 90 0.5 2.175
+ 90 0.5 2.2
+ 90 0.5 2.225
+ 90 0.5 2.25
+ 90 0.5 2.275
+ 90 0.5 2.3
+ 90 0.5 2.325
+ 90 0.5 2.35
+ 90 0.5 2.375
+ 90 0.5 2.4
+ 90 0.5 2.425
+ 90 0.5 2.45
+ 90 0.5 2.475
+ 90 0.5 2.5
+ 92 0.5 1.25
+ 92 0.5 1.275
+ 92 0.5 1.3
+ 92 0.5 1.325
+ 92 0.5 1.35
+ 92 0.5 1.375
+ 92 0.5 1.4
+ 92 0.5 1.425
+ 92 0.5 1.45
+ 92 0.5 1.475
+ 92 0.5 1.5
+ 92 0.5 1.525
+ 92 0.5 1.55
+ 92 0.5 1.575
+ 92 0.5 1.6
+ 92 0.5 1.625
+ 92 0.5 1.65
+ 92 0.5 1.675
+ 92 0.5 1.7
+ 92 0.5 1.725
+ 92 0.5 1.75
+ 92 0.5 1.775
+ 92 0.5 1.8
+ 92 0.5 1.825
+ 92 0.5 1.85
+ 92 0.5 1.875
+ 92 0.5 1.9
+ 92 0.5 1.925
+ 92 0.5 1.95
+ 92 0.5 1.975
+ 92 0.5 2.0
+ 92 0.5 2.025
+ 92 0.5 2.05
+ 92 0.5 2.075
+ 92 0.5 2.1
+ 92 0.5 2.125
+ 92 0.5 2.15
+ 92 0.5 2.175
+ 92 0.5 2.2
+ 92 0.5 2.225
+ 92 0.5 2.25
+ 92 0.5 2.275
+ 92 0.5 2.3
+ 92 0.5 2.325
+ 92 0.5 2.35
+ 92 0.5 2.375
+ 92 0.5 2.4
+ 92 0.5 2.425
+ 92 0.5 2.45
+ 92 0.5 2.475
+ 92 0.5 2.5
+ 94 0.5 1.25
+ 94 0.5 1.275
+ 94 0.5 1.3
+ 94 0.5 1.325
+ 94 0.5 1.35
+ 94 0.5 1.375
+ 94 0.5 1.4
+ 94 0.5 1.425
+ 94 0.5 1.45
+ 94 0.5 1.475
+ 94 0.5 1.5
+ 94 0.5 1.525
+ 94 0.5 1.55
+ 94 0.5 1.575
+ 94 0.5 1.6
+ 94 0.5 1.625
+ 94 0.5 1.65
+ 94 0.5 1.675
+ 94 0.5 1.7
+ 94 0.5 1.725
+ 94 0.5 1.75
+ 94 0.5 1.775
+ 94 0.5 1.8
+ 94 0.5 1.825
+ 94 0.5 1.85
+ 94 0.5 1.875
+ 94 0.5 1.9
+ 94 0.5 1.925
+ 94 0.5 1.95
+ 94 0.5 1.975
+ 94 0.5 2.0
+ 94 0.5 2.025
+ 94 0.5 2.05
+ 94 0.5 2.075
+ 94 0.5 2.1
+ 94 0.5 2.125
+ 94 0.5 2.15
+ 94 0.5 2.175
+ 94 0.5 2.2
+ 94 0.5 2.225
+ 94 0.5 2.25
+ 94 0.5 2.275
+ 94 0.5 2.3
+ 94 0.5 2.325
+ 94 0.5 2.35
+ 94 0.5 2.375
+ 94 0.5 2.4
+ 94 0.5 2.425
+ 94 0.5 2.45
+ 94 0.5 2.475
+ 94 0.5 2.5
+ 96 0.5 1.25
+ 96 0.5 1.275
+ 96 0.5 1.3
+ 96 0.5 1.325
+ 96 0.5 1.35
+ 96 0.5 1.375
+ 96 0.5 1.4
+ 96 0.5 1.425
+ 96 0.5 1.45
+ 96 0.5 1.475
+ 96 0.5 1.5
+ 96 0.5 1.525
+ 96 0.5 1.55
+ 96 0.5 1.575
+ 96 0.5 1.6
+ 96 0.5 1.625
+ 96 0.5 1.65
+ 96 0.5 1.675
+ 96 0.5 1.7
+ 96 0.5 1.725
+ 96 0.5 1.75
+ 96 0.5 1.775
+ 96 0.5 1.8
+ 96 0.5 1.825
+ 96 0.5 1.85
+ 96 0.5 1.875
+ 96 0.5 1.9
+ 96 0.5 1.925
+ 96 0.5 1.95
+ 96 0.5 1.975
+ 96 0.5 2.0
+ 96 0.5 2.025
+ 96 0.5 2.05
+ 96 0.5 2.075
+ 96 0.5 2.1
+ 96 0.5 2.125
+ 96 0.5 2.15
+ 96 0.5 2.175
+ 96 0.5 2.2
+ 96 0.5 2.225
+ 96 0.5 2.25
+ 96 0.5 2.275
+ 96 0.5 2.3
+ 96 0.5 2.325
+ 96 0.5 2.35
+ 96 0.5 2.375
+ 96 0.5 2.4
+ 96 0.5 2.425
+ 96 0.5 2.45
+ 96 0.5 2.475
+ 96 0.5 2.5
+ 98 0.5 1.25
+ 98 0.5 1.275
+ 98 0.5 1.3
+ 98 0.5 1.325
+ 98 0.5 1.35
+ 98 0.5 1.375
+ 98 0.5 1.4
+ 98 0.5 1.425
+ 98 0.5 1.45
+ 98 0.5 1.475
+ 98 0.5 1.5
+ 98 0.5 1.525
+ 98 0.5 1.55
+ 98 0.5 1.575
+ 98 0.5 1.6
+ 98 0.5 1.625
+ 98 0.5 1.65
+ 98 0.5 1.675
+ 98 0.5 1.7
+ 98 0.5 1.725
+ 98 0.5 1.75
+ 98 0.5 1.775
+ 98 0.5 1.8
+ 98 0.5 1.825
+ 98 0.5 1.85
+ 98 0.5 1.875
+ 98 0.5 1.9
+ 98 0.5 1.925
+ 98 0.5 1.95
+ 98 0.5 1.975
+ 98 0.5 2.0
+ 98 0.5 2.025
+ 98 0.5 2.05
+ 98 0.5 2.075
+ 98 0.5 2.1
+ 98 0.5 2.125
+ 98 0.5 2.15
+ 98 0.5 2.175
+ 98 0.5 2.2
+ 98 0.5 2.225
+ 98 0.5 2.25
+ 98 0.5 2.275
+ 98 0.5 2.3
+ 98 0.5 2.325
+ 98 0.5 2.35
+ 98 0.5 2.375
+ 98 0.5 2.4
+ 98 0.5 2.425
+ 98 0.5 2.45
+ 98 0.5 2.475
+ 98 0.5 2.5
+ 100 0.5 1.25
+ 100 0.5 1.275
+ 100 0.5 1.3
+ 100 0.5 1.325
+ 100 0.5 1.35
+ 100 0.5 1.375
+ 100 0.5 1.4
+ 100 0.5 1.425
+ 100 0.5 1.45
+ 100 0.5 1.475
+ 100 0.5 1.5
+ 100 0.5 1.525
+ 100 0.5 1.55
+ 100 0.5 1.575
+ 100 0.5 1.6
+ 100 0.5 1.625
+ 100 0.5 1.65
+ 100 0.5 1.675
+ 100 0.5 1.7
+ 100 0.5 1.725
+ 100 0.5 1.75
+ 100 0.5 1.775
+ 100 0.5 1.8
+ 100 0.5 1.825
+ 100 0.5 1.85
+ 100 0.5 1.875
+ 100 0.5 1.9
+ 100 0.5 1.925
+ 100 0.5 1.95
+ 100 0.5 1.975
+ 100 0.5 2.0
+ 100 0.5 2.025
+ 100 0.5 2.05
+ 100 0.5 2.075
+ 100 0.5 2.1
+ 100 0.5 2.125
+ 100 0.5 2.15
+ 100 0.5 2.175
+ 100 0.5 2.2
+ 100 0.5 2.225
+ 100 0.5 2.25
+ 100 0.5 2.275
+ 100 0.5 2.3
+ 100 0.5 2.325
+ 100 0.5 2.35
+ 100 0.5 2.375
+ 100 0.5 2.4
+ 100 0.5 2.425
+ 100 0.5 2.45
+ 100 0.5 2.475
+ 100 0.5 2.5
+ 0 0.6 1.25
+ 0 0.6 1.275
+ 0 0.6 1.3
+ 0 0.6 1.325
+ 0 0.6 1.35
+ 0 0.6 1.375
+ 0 0.6 1.4
+ 0 0.6 1.425
+ 0 0.6 1.45
+ 0 0.6 1.475
+ 0 0.6 1.5
+ 0 0.6 1.525
+ 0 0.6 1.55
+ 0 0.6 1.575
+ 0 0.6 1.6
+ 0 0.6 1.625
+ 0 0.6 1.65
+ 0 0.6 1.675
+ 0 0.6 1.7
+ 0 0.6 1.725
+ 0 0.6 1.75
+ 0 0.6 1.775
+ 0 0.6 1.8
+ 0 0.6 1.825
+ 0 0.6 1.85
+ 0 0.6 1.875
+ 0 0.6 1.9
+ 0 0.6 1.925
+ 0 0.6 1.95
+ 0 0.6 1.975
+ 0 0.6 2.0
+ 0 0.6 2.025
+ 0 0.6 2.05
+ 0 0.6 2.075
+ 0 0.6 2.1
+ 0 0.6 2.125
+ 0 0.6 2.15
+ 0 0.6 2.175
+ 0 0.6 2.2
+ 0 0.6 2.225
+ 0 0.6 2.25
+ 0 0.6 2.275
+ 0 0.6 2.3
+ 0 0.6 2.325
+ 0 0.6 2.35
+ 0 0.6 2.375
+ 0 0.6 2.4
+ 0 0.6 2.425
+ 0 0.6 2.45
+ 0 0.6 2.475
+ 0 0.6 2.5
+ 2 0.6 1.25
+ 2 0.6 1.275
+ 2 0.6 1.3
+ 2 0.6 1.325
+ 2 0.6 1.35
+ 2 0.6 1.375
+ 2 0.6 1.4
+ 2 0.6 1.425
+ 2 0.6 1.45
+ 2 0.6 1.475
+ 2 0.6 1.5
+ 2 0.6 1.525
+ 2 0.6 1.55
+ 2 0.6 1.575
+ 2 0.6 1.6
+ 2 0.6 1.625
+ 2 0.6 1.65
+ 2 0.6 1.675
+ 2 0.6 1.7
+ 2 0.6 1.725
+ 2 0.6 1.75
+ 2 0.6 1.775
+ 2 0.6 1.8
+ 2 0.6 1.825
+ 2 0.6 1.85
+ 2 0.6 1.875
+ 2 0.6 1.9
+ 2 0.6 1.925
+ 2 0.6 1.95
+ 2 0.6 1.975
+ 2 0.6 2.0
+ 2 0.6 2.025
+ 2 0.6 2.05
+ 2 0.6 2.075
+ 2 0.6 2.1
+ 2 0.6 2.125
+ 2 0.6 2.15
+ 2 0.6 2.175
+ 2 0.6 2.2
+ 2 0.6 2.225
+ 2 0.6 2.25
+ 2 0.6 2.275
+ 2 0.6 2.3
+ 2 0.6 2.325
+ 2 0.6 2.35
+ 2 0.6 2.375
+ 2 0.6 2.4
+ 2 0.6 2.425
+ 2 0.6 2.45
+ 2 0.6 2.475
+ 2 0.6 2.5
+ 4 0.6 1.25
+ 4 0.6 1.275
+ 4 0.6 1.3
+ 4 0.6 1.325
+ 4 0.6 1.35
+ 4 0.6 1.375
+ 4 0.6 1.4
+ 4 0.6 1.425
+ 4 0.6 1.45
+ 4 0.6 1.475
+ 4 0.6 1.5
+ 4 0.6 1.525
+ 4 0.6 1.55
+ 4 0.6 1.575
+ 4 0.6 1.6
+ 4 0.6 1.625
+ 4 0.6 1.65
+ 4 0.6 1.675
+ 4 0.6 1.7
+ 4 0.6 1.725
+ 4 0.6 1.75
+ 4 0.6 1.775
+ 4 0.6 1.8
+ 4 0.6 1.825
+ 4 0.6 1.85
+ 4 0.6 1.875
+ 4 0.6 1.9
+ 4 0.6 1.925
+ 4 0.6 1.95
+ 4 0.6 1.975
+ 4 0.6 2.0
+ 4 0.6 2.025
+ 4 0.6 2.05
+ 4 0.6 2.075
+ 4 0.6 2.1
+ 4 0.6 2.125
+ 4 0.6 2.15
+ 4 0.6 2.175
+ 4 0.6 2.2
+ 4 0.6 2.225
+ 4 0.6 2.25
+ 4 0.6 2.275
+ 4 0.6 2.3
+ 4 0.6 2.325
+ 4 0.6 2.35
+ 4 0.6 2.375
+ 4 0.6 2.4
+ 4 0.6 2.425
+ 4 0.6 2.45
+ 4 0.6 2.475
+ 4 0.6 2.5
+ 6 0.6 1.25
+ 6 0.6 1.275
+ 6 0.6 1.3
+ 6 0.6 1.325
+ 6 0.6 1.35
+ 6 0.6 1.375
+ 6 0.6 1.4
+ 6 0.6 1.425
+ 6 0.6 1.45
+ 6 0.6 1.475
+ 6 0.6 1.5
+ 6 0.6 1.525
+ 6 0.6 1.55
+ 6 0.6 1.575
+ 6 0.6 1.6
+ 6 0.6 1.625
+ 6 0.6 1.65
+ 6 0.6 1.675
+ 6 0.6 1.7
+ 6 0.6 1.725
+ 6 0.6 1.75
+ 6 0.6 1.775
+ 6 0.6 1.8
+ 6 0.6 1.825
+ 6 0.6 1.85
+ 6 0.6 1.875
+ 6 0.6 1.9
+ 6 0.6 1.925
+ 6 0.6 1.95
+ 6 0.6 1.975
+ 6 0.6 2.0
+ 6 0.6 2.025
+ 6 0.6 2.05
+ 6 0.6 2.075
+ 6 0.6 2.1
+ 6 0.6 2.125
+ 6 0.6 2.15
+ 6 0.6 2.175
+ 6 0.6 2.2
+ 6 0.6 2.225
+ 6 0.6 2.25
+ 6 0.6 2.275
+ 6 0.6 2.3
+ 6 0.6 2.325
+ 6 0.6 2.35
+ 6 0.6 2.375
+ 6 0.6 2.4
+ 6 0.6 2.425
+ 6 0.6 2.45
+ 6 0.6 2.475
+ 6 0.6 2.5
+ 8 0.6 1.25
+ 8 0.6 1.275
+ 8 0.6 1.3
+ 8 0.6 1.325
+ 8 0.6 1.35
+ 8 0.6 1.375
+ 8 0.6 1.4
+ 8 0.6 1.425
+ 8 0.6 1.45
+ 8 0.6 1.475
+ 8 0.6 1.5
+ 8 0.6 1.525
+ 8 0.6 1.55
+ 8 0.6 1.575
+ 8 0.6 1.6
+ 8 0.6 1.625
+ 8 0.6 1.65
+ 8 0.6 1.675
+ 8 0.6 1.7
+ 8 0.6 1.725
+ 8 0.6 1.75
+ 8 0.6 1.775
+ 8 0.6 1.8
+ 8 0.6 1.825
+ 8 0.6 1.85
+ 8 0.6 1.875
+ 8 0.6 1.9
+ 8 0.6 1.925
+ 8 0.6 1.95
+ 8 0.6 1.975
+ 8 0.6 2.0
+ 8 0.6 2.025
+ 8 0.6 2.05
+ 8 0.6 2.075
+ 8 0.6 2.1
+ 8 0.6 2.125
+ 8 0.6 2.15
+ 8 0.6 2.175
+ 8 0.6 2.2
+ 8 0.6 2.225
+ 8 0.6 2.25
+ 8 0.6 2.275
+ 8 0.6 2.3
+ 8 0.6 2.325
+ 8 0.6 2.35
+ 8 0.6 2.375
+ 8 0.6 2.4
+ 8 0.6 2.425
+ 8 0.6 2.45
+ 8 0.6 2.475
+ 8 0.6 2.5
+ 10 0.6 1.25
+ 10 0.6 1.275
+ 10 0.6 1.3
+ 10 0.6 1.325
+ 10 0.6 1.35
+ 10 0.6 1.375
+ 10 0.6 1.4
+ 10 0.6 1.425
+ 10 0.6 1.45
+ 10 0.6 1.475
+ 10 0.6 1.5
+ 10 0.6 1.525
+ 10 0.6 1.55
+ 10 0.6 1.575
+ 10 0.6 1.6
+ 10 0.6 1.625
+ 10 0.6 1.65
+ 10 0.6 1.675
+ 10 0.6 1.7
+ 10 0.6 1.725
+ 10 0.6 1.75
+ 10 0.6 1.775
+ 10 0.6 1.8
+ 10 0.6 1.825
+ 10 0.6 1.85
+ 10 0.6 1.875
+ 10 0.6 1.9
+ 10 0.6 1.925
+ 10 0.6 1.95
+ 10 0.6 1.975
+ 10 0.6 2.0
+ 10 0.6 2.025
+ 10 0.6 2.05
+ 10 0.6 2.075
+ 10 0.6 2.1
+ 10 0.6 2.125
+ 10 0.6 2.15
+ 10 0.6 2.175
+ 10 0.6 2.2
+ 10 0.6 2.225
+ 10 0.6 2.25
+ 10 0.6 2.275
+ 10 0.6 2.3
+ 10 0.6 2.325
+ 10 0.6 2.35
+ 10 0.6 2.375
+ 10 0.6 2.4
+ 10 0.6 2.425
+ 10 0.6 2.45
+ 10 0.6 2.475
+ 10 0.6 2.5
+ 12 0.6 1.25
+ 12 0.6 1.275
+ 12 0.6 1.3
+ 12 0.6 1.325
+ 12 0.6 1.35
+ 12 0.6 1.375
+ 12 0.6 1.4
+ 12 0.6 1.425
+ 12 0.6 1.45
+ 12 0.6 1.475
+ 12 0.6 1.5
+ 12 0.6 1.525
+ 12 0.6 1.55
+ 12 0.6 1.575
+ 12 0.6 1.6
+ 12 0.6 1.625
+ 12 0.6 1.65
+ 12 0.6 1.675
+ 12 0.6 1.7
+ 12 0.6 1.725
+ 12 0.6 1.75
+ 12 0.6 1.775
+ 12 0.6 1.8
+ 12 0.6 1.825
+ 12 0.6 1.85
+ 12 0.6 1.875
+ 12 0.6 1.9
+ 12 0.6 1.925
+ 12 0.6 1.95
+ 12 0.6 1.975
+ 12 0.6 2.0
+ 12 0.6 2.025
+ 12 0.6 2.05
+ 12 0.6 2.075
+ 12 0.6 2.1
+ 12 0.6 2.125
+ 12 0.6 2.15
+ 12 0.6 2.175
+ 12 0.6 2.2
+ 12 0.6 2.225
+ 12 0.6 2.25
+ 12 0.6 2.275
+ 12 0.6 2.3
+ 12 0.6 2.325
+ 12 0.6 2.35
+ 12 0.6 2.375
+ 12 0.6 2.4
+ 12 0.6 2.425
+ 12 0.6 2.45
+ 12 0.6 2.475
+ 12 0.6 2.5
+ 14 0.6 1.25
+ 14 0.6 1.275
+ 14 0.6 1.3
+ 14 0.6 1.325
+ 14 0.6 1.35
+ 14 0.6 1.375
+ 14 0.6 1.4
+ 14 0.6 1.425
+ 14 0.6 1.45
+ 14 0.6 1.475
+ 14 0.6 1.5
+ 14 0.6 1.525
+ 14 0.6 1.55
+ 14 0.6 1.575
+ 14 0.6 1.6
+ 14 0.6 1.625
+ 14 0.6 1.65
+ 14 0.6 1.675
+ 14 0.6 1.7
+ 14 0.6 1.725
+ 14 0.6 1.75
+ 14 0.6 1.775
+ 14 0.6 1.8
+ 14 0.6 1.825
+ 14 0.6 1.85
+ 14 0.6 1.875
+ 14 0.6 1.9
+ 14 0.6 1.925
+ 14 0.6 1.95
+ 14 0.6 1.975
+ 14 0.6 2.0
+ 14 0.6 2.025
+ 14 0.6 2.05
+ 14 0.6 2.075
+ 14 0.6 2.1
+ 14 0.6 2.125
+ 14 0.6 2.15
+ 14 0.6 2.175
+ 14 0.6 2.2
+ 14 0.6 2.225
+ 14 0.6 2.25
+ 14 0.6 2.275
+ 14 0.6 2.3
+ 14 0.6 2.325
+ 14 0.6 2.35
+ 14 0.6 2.375
+ 14 0.6 2.4
+ 14 0.6 2.425
+ 14 0.6 2.45
+ 14 0.6 2.475
+ 14 0.6 2.5
+ 16 0.6 1.25
+ 16 0.6 1.275
+ 16 0.6 1.3
+ 16 0.6 1.325
+ 16 0.6 1.35
+ 16 0.6 1.375
+ 16 0.6 1.4
+ 16 0.6 1.425
+ 16 0.6 1.45
+ 16 0.6 1.475
+ 16 0.6 1.5
+ 16 0.6 1.525
+ 16 0.6 1.55
+ 16 0.6 1.575
+ 16 0.6 1.6
+ 16 0.6 1.625
+ 16 0.6 1.65
+ 16 0.6 1.675
+ 16 0.6 1.7
+ 16 0.6 1.725
+ 16 0.6 1.75
+ 16 0.6 1.775
+ 16 0.6 1.8
+ 16 0.6 1.825
+ 16 0.6 1.85
+ 16 0.6 1.875
+ 16 0.6 1.9
+ 16 0.6 1.925
+ 16 0.6 1.95
+ 16 0.6 1.975
+ 16 0.6 2.0
+ 16 0.6 2.025
+ 16 0.6 2.05
+ 16 0.6 2.075
+ 16 0.6 2.1
+ 16 0.6 2.125
+ 16 0.6 2.15
+ 16 0.6 2.175
+ 16 0.6 2.2
+ 16 0.6 2.225
+ 16 0.6 2.25
+ 16 0.6 2.275
+ 16 0.6 2.3
+ 16 0.6 2.325
+ 16 0.6 2.35
+ 16 0.6 2.375
+ 16 0.6 2.4
+ 16 0.6 2.425
+ 16 0.6 2.45
+ 16 0.6 2.475
+ 16 0.6 2.5
+ 18 0.6 1.25
+ 18 0.6 1.275
+ 18 0.6 1.3
+ 18 0.6 1.325
+ 18 0.6 1.35
+ 18 0.6 1.375
+ 18 0.6 1.4
+ 18 0.6 1.425
+ 18 0.6 1.45
+ 18 0.6 1.475
+ 18 0.6 1.5
+ 18 0.6 1.525
+ 18 0.6 1.55
+ 18 0.6 1.575
+ 18 0.6 1.6
+ 18 0.6 1.625
+ 18 0.6 1.65
+ 18 0.6 1.675
+ 18 0.6 1.7
+ 18 0.6 1.725
+ 18 0.6 1.75
+ 18 0.6 1.775
+ 18 0.6 1.8
+ 18 0.6 1.825
+ 18 0.6 1.85
+ 18 0.6 1.875
+ 18 0.6 1.9
+ 18 0.6 1.925
+ 18 0.6 1.95
+ 18 0.6 1.975
+ 18 0.6 2.0
+ 18 0.6 2.025
+ 18 0.6 2.05
+ 18 0.6 2.075
+ 18 0.6 2.1
+ 18 0.6 2.125
+ 18 0.6 2.15
+ 18 0.6 2.175
+ 18 0.6 2.2
+ 18 0.6 2.225
+ 18 0.6 2.25
+ 18 0.6 2.275
+ 18 0.6 2.3
+ 18 0.6 2.325
+ 18 0.6 2.35
+ 18 0.6 2.375
+ 18 0.6 2.4
+ 18 0.6 2.425
+ 18 0.6 2.45
+ 18 0.6 2.475
+ 18 0.6 2.5
+ 20 0.6 1.25
+ 20 0.6 1.275
+ 20 0.6 1.3
+ 20 0.6 1.325
+ 20 0.6 1.35
+ 20 0.6 1.375
+ 20 0.6 1.4
+ 20 0.6 1.425
+ 20 0.6 1.45
+ 20 0.6 1.475
+ 20 0.6 1.5
+ 20 0.6 1.525
+ 20 0.6 1.55
+ 20 0.6 1.575
+ 20 0.6 1.6
+ 20 0.6 1.625
+ 20 0.6 1.65
+ 20 0.6 1.675
+ 20 0.6 1.7
+ 20 0.6 1.725
+ 20 0.6 1.75
+ 20 0.6 1.775
+ 20 0.6 1.8
+ 20 0.6 1.825
+ 20 0.6 1.85
+ 20 0.6 1.875
+ 20 0.6 1.9
+ 20 0.6 1.925
+ 20 0.6 1.95
+ 20 0.6 1.975
+ 20 0.6 2.0
+ 20 0.6 2.025
+ 20 0.6 2.05
+ 20 0.6 2.075
+ 20 0.6 2.1
+ 20 0.6 2.125
+ 20 0.6 2.15
+ 20 0.6 2.175
+ 20 0.6 2.2
+ 20 0.6 2.225
+ 20 0.6 2.25
+ 20 0.6 2.275
+ 20 0.6 2.3
+ 20 0.6 2.325
+ 20 0.6 2.35
+ 20 0.6 2.375
+ 20 0.6 2.4
+ 20 0.6 2.425
+ 20 0.6 2.45
+ 20 0.6 2.475
+ 20 0.6 2.5
+ 22 0.6 1.25
+ 22 0.6 1.275
+ 22 0.6 1.3
+ 22 0.6 1.325
+ 22 0.6 1.35
+ 22 0.6 1.375
+ 22 0.6 1.4
+ 22 0.6 1.425
+ 22 0.6 1.45
+ 22 0.6 1.475
+ 22 0.6 1.5
+ 22 0.6 1.525
+ 22 0.6 1.55
+ 22 0.6 1.575
+ 22 0.6 1.6
+ 22 0.6 1.625
+ 22 0.6 1.65
+ 22 0.6 1.675
+ 22 0.6 1.7
+ 22 0.6 1.725
+ 22 0.6 1.75
+ 22 0.6 1.775
+ 22 0.6 1.8
+ 22 0.6 1.825
+ 22 0.6 1.85
+ 22 0.6 1.875
+ 22 0.6 1.9
+ 22 0.6 1.925
+ 22 0.6 1.95
+ 22 0.6 1.975
+ 22 0.6 2.0
+ 22 0.6 2.025
+ 22 0.6 2.05
+ 22 0.6 2.075
+ 22 0.6 2.1
+ 22 0.6 2.125
+ 22 0.6 2.15
+ 22 0.6 2.175
+ 22 0.6 2.2
+ 22 0.6 2.225
+ 22 0.6 2.25
+ 22 0.6 2.275
+ 22 0.6 2.3
+ 22 0.6 2.325
+ 22 0.6 2.35
+ 22 0.6 2.375
+ 22 0.6 2.4
+ 22 0.6 2.425
+ 22 0.6 2.45
+ 22 0.6 2.475
+ 22 0.6 2.5
+ 24 0.6 1.25
+ 24 0.6 1.275
+ 24 0.6 1.3
+ 24 0.6 1.325
+ 24 0.6 1.35
+ 24 0.6 1.375
+ 24 0.6 1.4
+ 24 0.6 1.425
+ 24 0.6 1.45
+ 24 0.6 1.475
+ 24 0.6 1.5
+ 24 0.6 1.525
+ 24 0.6 1.55
+ 24 0.6 1.575
+ 24 0.6 1.6
+ 24 0.6 1.625
+ 24 0.6 1.65
+ 24 0.6 1.675
+ 24 0.6 1.7
+ 24 0.6 1.725
+ 24 0.6 1.75
+ 24 0.6 1.775
+ 24 0.6 1.8
+ 24 0.6 1.825
+ 24 0.6 1.85
+ 24 0.6 1.875
+ 24 0.6 1.9
+ 24 0.6 1.925
+ 24 0.6 1.95
+ 24 0.6 1.975
+ 24 0.6 2.0
+ 24 0.6 2.025
+ 24 0.6 2.05
+ 24 0.6 2.075
+ 24 0.6 2.1
+ 24 0.6 2.125
+ 24 0.6 2.15
+ 24 0.6 2.175
+ 24 0.6 2.2
+ 24 0.6 2.225
+ 24 0.6 2.25
+ 24 0.6 2.275
+ 24 0.6 2.3
+ 24 0.6 2.325
+ 24 0.6 2.35
+ 24 0.6 2.375
+ 24 0.6 2.4
+ 24 0.6 2.425
+ 24 0.6 2.45
+ 24 0.6 2.475
+ 24 0.6 2.5
+ 26 0.6 1.25
+ 26 0.6 1.275
+ 26 0.6 1.3
+ 26 0.6 1.325
+ 26 0.6 1.35
+ 26 0.6 1.375
+ 26 0.6 1.4
+ 26 0.6 1.425
+ 26 0.6 1.45
+ 26 0.6 1.475
+ 26 0.6 1.5
+ 26 0.6 1.525
+ 26 0.6 1.55
+ 26 0.6 1.575
+ 26 0.6 1.6
+ 26 0.6 1.625
+ 26 0.6 1.65
+ 26 0.6 1.675
+ 26 0.6 1.7
+ 26 0.6 1.725
+ 26 0.6 1.75
+ 26 0.6 1.775
+ 26 0.6 1.8
+ 26 0.6 1.825
+ 26 0.6 1.85
+ 26 0.6 1.875
+ 26 0.6 1.9
+ 26 0.6 1.925
+ 26 0.6 1.95
+ 26 0.6 1.975
+ 26 0.6 2.0
+ 26 0.6 2.025
+ 26 0.6 2.05
+ 26 0.6 2.075
+ 26 0.6 2.1
+ 26 0.6 2.125
+ 26 0.6 2.15
+ 26 0.6 2.175
+ 26 0.6 2.2
+ 26 0.6 2.225
+ 26 0.6 2.25
+ 26 0.6 2.275
+ 26 0.6 2.3
+ 26 0.6 2.325
+ 26 0.6 2.35
+ 26 0.6 2.375
+ 26 0.6 2.4
+ 26 0.6 2.425
+ 26 0.6 2.45
+ 26 0.6 2.475
+ 26 0.6 2.5
+ 28 0.6 1.25
+ 28 0.6 1.275
+ 28 0.6 1.3
+ 28 0.6 1.325
+ 28 0.6 1.35
+ 28 0.6 1.375
+ 28 0.6 1.4
+ 28 0.6 1.425
+ 28 0.6 1.45
+ 28 0.6 1.475
+ 28 0.6 1.5
+ 28 0.6 1.525
+ 28 0.6 1.55
+ 28 0.6 1.575
+ 28 0.6 1.6
+ 28 0.6 1.625
+ 28 0.6 1.65
+ 28 0.6 1.675
+ 28 0.6 1.7
+ 28 0.6 1.725
+ 28 0.6 1.75
+ 28 0.6 1.775
+ 28 0.6 1.8
+ 28 0.6 1.825
+ 28 0.6 1.85
+ 28 0.6 1.875
+ 28 0.6 1.9
+ 28 0.6 1.925
+ 28 0.6 1.95
+ 28 0.6 1.975
+ 28 0.6 2.0
+ 28 0.6 2.025
+ 28 0.6 2.05
+ 28 0.6 2.075
+ 28 0.6 2.1
+ 28 0.6 2.125
+ 28 0.6 2.15
+ 28 0.6 2.175
+ 28 0.6 2.2
+ 28 0.6 2.225
+ 28 0.6 2.25
+ 28 0.6 2.275
+ 28 0.6 2.3
+ 28 0.6 2.325
+ 28 0.6 2.35
+ 28 0.6 2.375
+ 28 0.6 2.4
+ 28 0.6 2.425
+ 28 0.6 2.45
+ 28 0.6 2.475
+ 28 0.6 2.5
+ 30 0.6 1.25
+ 30 0.6 1.275
+ 30 0.6 1.3
+ 30 0.6 1.325
+ 30 0.6 1.35
+ 30 0.6 1.375
+ 30 0.6 1.4
+ 30 0.6 1.425
+ 30 0.6 1.45
+ 30 0.6 1.475
+ 30 0.6 1.5
+ 30 0.6 1.525
+ 30 0.6 1.55
+ 30 0.6 1.575
+ 30 0.6 1.6
+ 30 0.6 1.625
+ 30 0.6 1.65
+ 30 0.6 1.675
+ 30 0.6 1.7
+ 30 0.6 1.725
+ 30 0.6 1.75
+ 30 0.6 1.775
+ 30 0.6 1.8
+ 30 0.6 1.825
+ 30 0.6 1.85
+ 30 0.6 1.875
+ 30 0.6 1.9
+ 30 0.6 1.925
+ 30 0.6 1.95
+ 30 0.6 1.975
+ 30 0.6 2.0
+ 30 0.6 2.025
+ 30 0.6 2.05
+ 30 0.6 2.075
+ 30 0.6 2.1
+ 30 0.6 2.125
+ 30 0.6 2.15
+ 30 0.6 2.175
+ 30 0.6 2.2
+ 30 0.6 2.225
+ 30 0.6 2.25
+ 30 0.6 2.275
+ 30 0.6 2.3
+ 30 0.6 2.325
+ 30 0.6 2.35
+ 30 0.6 2.375
+ 30 0.6 2.4
+ 30 0.6 2.425
+ 30 0.6 2.45
+ 30 0.6 2.475
+ 30 0.6 2.5
+ 32 0.6 1.25
+ 32 0.6 1.275
+ 32 0.6 1.3
+ 32 0.6 1.325
+ 32 0.6 1.35
+ 32 0.6 1.375
+ 32 0.6 1.4
+ 32 0.6 1.425
+ 32 0.6 1.45
+ 32 0.6 1.475
+ 32 0.6 1.5
+ 32 0.6 1.525
+ 32 0.6 1.55
+ 32 0.6 1.575
+ 32 0.6 1.6
+ 32 0.6 1.625
+ 32 0.6 1.65
+ 32 0.6 1.675
+ 32 0.6 1.7
+ 32 0.6 1.725
+ 32 0.6 1.75
+ 32 0.6 1.775
+ 32 0.6 1.8
+ 32 0.6 1.825
+ 32 0.6 1.85
+ 32 0.6 1.875
+ 32 0.6 1.9
+ 32 0.6 1.925
+ 32 0.6 1.95
+ 32 0.6 1.975
+ 32 0.6 2.0
+ 32 0.6 2.025
+ 32 0.6 2.05
+ 32 0.6 2.075
+ 32 0.6 2.1
+ 32 0.6 2.125
+ 32 0.6 2.15
+ 32 0.6 2.175
+ 32 0.6 2.2
+ 32 0.6 2.225
+ 32 0.6 2.25
+ 32 0.6 2.275
+ 32 0.6 2.3
+ 32 0.6 2.325
+ 32 0.6 2.35
+ 32 0.6 2.375
+ 32 0.6 2.4
+ 32 0.6 2.425
+ 32 0.6 2.45
+ 32 0.6 2.475
+ 32 0.6 2.5
+ 34 0.6 1.25
+ 34 0.6 1.275
+ 34 0.6 1.3
+ 34 0.6 1.325
+ 34 0.6 1.35
+ 34 0.6 1.375
+ 34 0.6 1.4
+ 34 0.6 1.425
+ 34 0.6 1.45
+ 34 0.6 1.475
+ 34 0.6 1.5
+ 34 0.6 1.525
+ 34 0.6 1.55
+ 34 0.6 1.575
+ 34 0.6 1.6
+ 34 0.6 1.625
+ 34 0.6 1.65
+ 34 0.6 1.675
+ 34 0.6 1.7
+ 34 0.6 1.725
+ 34 0.6 1.75
+ 34 0.6 1.775
+ 34 0.6 1.8
+ 34 0.6 1.825
+ 34 0.6 1.85
+ 34 0.6 1.875
+ 34 0.6 1.9
+ 34 0.6 1.925
+ 34 0.6 1.95
+ 34 0.6 1.975
+ 34 0.6 2.0
+ 34 0.6 2.025
+ 34 0.6 2.05
+ 34 0.6 2.075
+ 34 0.6 2.1
+ 34 0.6 2.125
+ 34 0.6 2.15
+ 34 0.6 2.175
+ 34 0.6 2.2
+ 34 0.6 2.225
+ 34 0.6 2.25
+ 34 0.6 2.275
+ 34 0.6 2.3
+ 34 0.6 2.325
+ 34 0.6 2.35
+ 34 0.6 2.375
+ 34 0.6 2.4
+ 34 0.6 2.425
+ 34 0.6 2.45
+ 34 0.6 2.475
+ 34 0.6 2.5
+ 36 0.6 1.25
+ 36 0.6 1.275
+ 36 0.6 1.3
+ 36 0.6 1.325
+ 36 0.6 1.35
+ 36 0.6 1.375
+ 36 0.6 1.4
+ 36 0.6 1.425
+ 36 0.6 1.45
+ 36 0.6 1.475
+ 36 0.6 1.5
+ 36 0.6 1.525
+ 36 0.6 1.55
+ 36 0.6 1.575
+ 36 0.6 1.6
+ 36 0.6 1.625
+ 36 0.6 1.65
+ 36 0.6 1.675
+ 36 0.6 1.7
+ 36 0.6 1.725
+ 36 0.6 1.75
+ 36 0.6 1.775
+ 36 0.6 1.8
+ 36 0.6 1.825
+ 36 0.6 1.85
+ 36 0.6 1.875
+ 36 0.6 1.9
+ 36 0.6 1.925
+ 36 0.6 1.95
+ 36 0.6 1.975
+ 36 0.6 2.0
+ 36 0.6 2.025
+ 36 0.6 2.05
+ 36 0.6 2.075
+ 36 0.6 2.1
+ 36 0.6 2.125
+ 36 0.6 2.15
+ 36 0.6 2.175
+ 36 0.6 2.2
+ 36 0.6 2.225
+ 36 0.6 2.25
+ 36 0.6 2.275
+ 36 0.6 2.3
+ 36 0.6 2.325
+ 36 0.6 2.35
+ 36 0.6 2.375
+ 36 0.6 2.4
+ 36 0.6 2.425
+ 36 0.6 2.45
+ 36 0.6 2.475
+ 36 0.6 2.5
+ 38 0.6 1.25
+ 38 0.6 1.275
+ 38 0.6 1.3
+ 38 0.6 1.325
+ 38 0.6 1.35
+ 38 0.6 1.375
+ 38 0.6 1.4
+ 38 0.6 1.425
+ 38 0.6 1.45
+ 38 0.6 1.475
+ 38 0.6 1.5
+ 38 0.6 1.525
+ 38 0.6 1.55
+ 38 0.6 1.575
+ 38 0.6 1.6
+ 38 0.6 1.625
+ 38 0.6 1.65
+ 38 0.6 1.675
+ 38 0.6 1.7
+ 38 0.6 1.725
+ 38 0.6 1.75
+ 38 0.6 1.775
+ 38 0.6 1.8
+ 38 0.6 1.825
+ 38 0.6 1.85
+ 38 0.6 1.875
+ 38 0.6 1.9
+ 38 0.6 1.925
+ 38 0.6 1.95
+ 38 0.6 1.975
+ 38 0.6 2.0
+ 38 0.6 2.025
+ 38 0.6 2.05
+ 38 0.6 2.075
+ 38 0.6 2.1
+ 38 0.6 2.125
+ 38 0.6 2.15
+ 38 0.6 2.175
+ 38 0.6 2.2
+ 38 0.6 2.225
+ 38 0.6 2.25
+ 38 0.6 2.275
+ 38 0.6 2.3
+ 38 0.6 2.325
+ 38 0.6 2.35
+ 38 0.6 2.375
+ 38 0.6 2.4
+ 38 0.6 2.425
+ 38 0.6 2.45
+ 38 0.6 2.475
+ 38 0.6 2.5
+ 40 0.6 1.25
+ 40 0.6 1.275
+ 40 0.6 1.3
+ 40 0.6 1.325
+ 40 0.6 1.35
+ 40 0.6 1.375
+ 40 0.6 1.4
+ 40 0.6 1.425
+ 40 0.6 1.45
+ 40 0.6 1.475
+ 40 0.6 1.5
+ 40 0.6 1.525
+ 40 0.6 1.55
+ 40 0.6 1.575
+ 40 0.6 1.6
+ 40 0.6 1.625
+ 40 0.6 1.65
+ 40 0.6 1.675
+ 40 0.6 1.7
+ 40 0.6 1.725
+ 40 0.6 1.75
+ 40 0.6 1.775
+ 40 0.6 1.8
+ 40 0.6 1.825
+ 40 0.6 1.85
+ 40 0.6 1.875
+ 40 0.6 1.9
+ 40 0.6 1.925
+ 40 0.6 1.95
+ 40 0.6 1.975
+ 40 0.6 2.0
+ 40 0.6 2.025
+ 40 0.6 2.05
+ 40 0.6 2.075
+ 40 0.6 2.1
+ 40 0.6 2.125
+ 40 0.6 2.15
+ 40 0.6 2.175
+ 40 0.6 2.2
+ 40 0.6 2.225
+ 40 0.6 2.25
+ 40 0.6 2.275
+ 40 0.6 2.3
+ 40 0.6 2.325
+ 40 0.6 2.35
+ 40 0.6 2.375
+ 40 0.6 2.4
+ 40 0.6 2.425
+ 40 0.6 2.45
+ 40 0.6 2.475
+ 40 0.6 2.5
+ 42 0.6 1.25
+ 42 0.6 1.275
+ 42 0.6 1.3
+ 42 0.6 1.325
+ 42 0.6 1.35
+ 42 0.6 1.375
+ 42 0.6 1.4
+ 42 0.6 1.425
+ 42 0.6 1.45
+ 42 0.6 1.475
+ 42 0.6 1.5
+ 42 0.6 1.525
+ 42 0.6 1.55
+ 42 0.6 1.575
+ 42 0.6 1.6
+ 42 0.6 1.625
+ 42 0.6 1.65
+ 42 0.6 1.675
+ 42 0.6 1.7
+ 42 0.6 1.725
+ 42 0.6 1.75
+ 42 0.6 1.775
+ 42 0.6 1.8
+ 42 0.6 1.825
+ 42 0.6 1.85
+ 42 0.6 1.875
+ 42 0.6 1.9
+ 42 0.6 1.925
+ 42 0.6 1.95
+ 42 0.6 1.975
+ 42 0.6 2.0
+ 42 0.6 2.025
+ 42 0.6 2.05
+ 42 0.6 2.075
+ 42 0.6 2.1
+ 42 0.6 2.125
+ 42 0.6 2.15
+ 42 0.6 2.175
+ 42 0.6 2.2
+ 42 0.6 2.225
+ 42 0.6 2.25
+ 42 0.6 2.275
+ 42 0.6 2.3
+ 42 0.6 2.325
+ 42 0.6 2.35
+ 42 0.6 2.375
+ 42 0.6 2.4
+ 42 0.6 2.425
+ 42 0.6 2.45
+ 42 0.6 2.475
+ 42 0.6 2.5
+ 44 0.6 1.25
+ 44 0.6 1.275
+ 44 0.6 1.3
+ 44 0.6 1.325
+ 44 0.6 1.35
+ 44 0.6 1.375
+ 44 0.6 1.4
+ 44 0.6 1.425
+ 44 0.6 1.45
+ 44 0.6 1.475
+ 44 0.6 1.5
+ 44 0.6 1.525
+ 44 0.6 1.55
+ 44 0.6 1.575
+ 44 0.6 1.6
+ 44 0.6 1.625
+ 44 0.6 1.65
+ 44 0.6 1.675
+ 44 0.6 1.7
+ 44 0.6 1.725
+ 44 0.6 1.75
+ 44 0.6 1.775
+ 44 0.6 1.8
+ 44 0.6 1.825
+ 44 0.6 1.85
+ 44 0.6 1.875
+ 44 0.6 1.9
+ 44 0.6 1.925
+ 44 0.6 1.95
+ 44 0.6 1.975
+ 44 0.6 2.0
+ 44 0.6 2.025
+ 44 0.6 2.05
+ 44 0.6 2.075
+ 44 0.6 2.1
+ 44 0.6 2.125
+ 44 0.6 2.15
+ 44 0.6 2.175
+ 44 0.6 2.2
+ 44 0.6 2.225
+ 44 0.6 2.25
+ 44 0.6 2.275
+ 44 0.6 2.3
+ 44 0.6 2.325
+ 44 0.6 2.35
+ 44 0.6 2.375
+ 44 0.6 2.4
+ 44 0.6 2.425
+ 44 0.6 2.45
+ 44 0.6 2.475
+ 44 0.6 2.5
+ 46 0.6 1.25
+ 46 0.6 1.275
+ 46 0.6 1.3
+ 46 0.6 1.325
+ 46 0.6 1.35
+ 46 0.6 1.375
+ 46 0.6 1.4
+ 46 0.6 1.425
+ 46 0.6 1.45
+ 46 0.6 1.475
+ 46 0.6 1.5
+ 46 0.6 1.525
+ 46 0.6 1.55
+ 46 0.6 1.575
+ 46 0.6 1.6
+ 46 0.6 1.625
+ 46 0.6 1.65
+ 46 0.6 1.675
+ 46 0.6 1.7
+ 46 0.6 1.725
+ 46 0.6 1.75
+ 46 0.6 1.775
+ 46 0.6 1.8
+ 46 0.6 1.825
+ 46 0.6 1.85
+ 46 0.6 1.875
+ 46 0.6 1.9
+ 46 0.6 1.925
+ 46 0.6 1.95
+ 46 0.6 1.975
+ 46 0.6 2.0
+ 46 0.6 2.025
+ 46 0.6 2.05
+ 46 0.6 2.075
+ 46 0.6 2.1
+ 46 0.6 2.125
+ 46 0.6 2.15
+ 46 0.6 2.175
+ 46 0.6 2.2
+ 46 0.6 2.225
+ 46 0.6 2.25
+ 46 0.6 2.275
+ 46 0.6 2.3
+ 46 0.6 2.325
+ 46 0.6 2.35
+ 46 0.6 2.375
+ 46 0.6 2.4
+ 46 0.6 2.425
+ 46 0.6 2.45
+ 46 0.6 2.475
+ 46 0.6 2.5
+ 48 0.6 1.25
+ 48 0.6 1.275
+ 48 0.6 1.3
+ 48 0.6 1.325
+ 48 0.6 1.35
+ 48 0.6 1.375
+ 48 0.6 1.4
+ 48 0.6 1.425
+ 48 0.6 1.45
+ 48 0.6 1.475
+ 48 0.6 1.5
+ 48 0.6 1.525
+ 48 0.6 1.55
+ 48 0.6 1.575
+ 48 0.6 1.6
+ 48 0.6 1.625
+ 48 0.6 1.65
+ 48 0.6 1.675
+ 48 0.6 1.7
+ 48 0.6 1.725
+ 48 0.6 1.75
+ 48 0.6 1.775
+ 48 0.6 1.8
+ 48 0.6 1.825
+ 48 0.6 1.85
+ 48 0.6 1.875
+ 48 0.6 1.9
+ 48 0.6 1.925
+ 48 0.6 1.95
+ 48 0.6 1.975
+ 48 0.6 2.0
+ 48 0.6 2.025
+ 48 0.6 2.05
+ 48 0.6 2.075
+ 48 0.6 2.1
+ 48 0.6 2.125
+ 48 0.6 2.15
+ 48 0.6 2.175
+ 48 0.6 2.2
+ 48 0.6 2.225
+ 48 0.6 2.25
+ 48 0.6 2.275
+ 48 0.6 2.3
+ 48 0.6 2.325
+ 48 0.6 2.35
+ 48 0.6 2.375
+ 48 0.6 2.4
+ 48 0.6 2.425
+ 48 0.6 2.45
+ 48 0.6 2.475
+ 48 0.6 2.5
+ 50 0.6 1.25
+ 50 0.6 1.275
+ 50 0.6 1.3
+ 50 0.6 1.325
+ 50 0.6 1.35
+ 50 0.6 1.375
+ 50 0.6 1.4
+ 50 0.6 1.425
+ 50 0.6 1.45
+ 50 0.6 1.475
+ 50 0.6 1.5
+ 50 0.6 1.525
+ 50 0.6 1.55
+ 50 0.6 1.575
+ 50 0.6 1.6
+ 50 0.6 1.625
+ 50 0.6 1.65
+ 50 0.6 1.675
+ 50 0.6 1.7
+ 50 0.6 1.725
+ 50 0.6 1.75
+ 50 0.6 1.775
+ 50 0.6 1.8
+ 50 0.6 1.825
+ 50 0.6 1.85
+ 50 0.6 1.875
+ 50 0.6 1.9
+ 50 0.6 1.925
+ 50 0.6 1.95
+ 50 0.6 1.975
+ 50 0.6 2.0
+ 50 0.6 2.025
+ 50 0.6 2.05
+ 50 0.6 2.075
+ 50 0.6 2.1
+ 50 0.6 2.125
+ 50 0.6 2.15
+ 50 0.6 2.175
+ 50 0.6 2.2
+ 50 0.6 2.225
+ 50 0.6 2.25
+ 50 0.6 2.275
+ 50 0.6 2.3
+ 50 0.6 2.325
+ 50 0.6 2.35
+ 50 0.6 2.375
+ 50 0.6 2.4
+ 50 0.6 2.425
+ 50 0.6 2.45
+ 50 0.6 2.475
+ 50 0.6 2.5
+ 52 0.6 1.25
+ 52 0.6 1.275
+ 52 0.6 1.3
+ 52 0.6 1.325
+ 52 0.6 1.35
+ 52 0.6 1.375
+ 52 0.6 1.4
+ 52 0.6 1.425
+ 52 0.6 1.45
+ 52 0.6 1.475
+ 52 0.6 1.5
+ 52 0.6 1.525
+ 52 0.6 1.55
+ 52 0.6 1.575
+ 52 0.6 1.6
+ 52 0.6 1.625
+ 52 0.6 1.65
+ 52 0.6 1.675
+ 52 0.6 1.7
+ 52 0.6 1.725
+ 52 0.6 1.75
+ 52 0.6 1.775
+ 52 0.6 1.8
+ 52 0.6 1.825
+ 52 0.6 1.85
+ 52 0.6 1.875
+ 52 0.6 1.9
+ 52 0.6 1.925
+ 52 0.6 1.95
+ 52 0.6 1.975
+ 52 0.6 2.0
+ 52 0.6 2.025
+ 52 0.6 2.05
+ 52 0.6 2.075
+ 52 0.6 2.1
+ 52 0.6 2.125
+ 52 0.6 2.15
+ 52 0.6 2.175
+ 52 0.6 2.2
+ 52 0.6 2.225
+ 52 0.6 2.25
+ 52 0.6 2.275
+ 52 0.6 2.3
+ 52 0.6 2.325
+ 52 0.6 2.35
+ 52 0.6 2.375
+ 52 0.6 2.4
+ 52 0.6 2.425
+ 52 0.6 2.45
+ 52 0.6 2.475
+ 52 0.6 2.5
+ 54 0.6 1.25
+ 54 0.6 1.275
+ 54 0.6 1.3
+ 54 0.6 1.325
+ 54 0.6 1.35
+ 54 0.6 1.375
+ 54 0.6 1.4
+ 54 0.6 1.425
+ 54 0.6 1.45
+ 54 0.6 1.475
+ 54 0.6 1.5
+ 54 0.6 1.525
+ 54 0.6 1.55
+ 54 0.6 1.575
+ 54 0.6 1.6
+ 54 0.6 1.625
+ 54 0.6 1.65
+ 54 0.6 1.675
+ 54 0.6 1.7
+ 54 0.6 1.725
+ 54 0.6 1.75
+ 54 0.6 1.775
+ 54 0.6 1.8
+ 54 0.6 1.825
+ 54 0.6 1.85
+ 54 0.6 1.875
+ 54 0.6 1.9
+ 54 0.6 1.925
+ 54 0.6 1.95
+ 54 0.6 1.975
+ 54 0.6 2.0
+ 54 0.6 2.025
+ 54 0.6 2.05
+ 54 0.6 2.075
+ 54 0.6 2.1
+ 54 0.6 2.125
+ 54 0.6 2.15
+ 54 0.6 2.175
+ 54 0.6 2.2
+ 54 0.6 2.225
+ 54 0.6 2.25
+ 54 0.6 2.275
+ 54 0.6 2.3
+ 54 0.6 2.325
+ 54 0.6 2.35
+ 54 0.6 2.375
+ 54 0.6 2.4
+ 54 0.6 2.425
+ 54 0.6 2.45
+ 54 0.6 2.475
+ 54 0.6 2.5
+ 56 0.6 1.25
+ 56 0.6 1.275
+ 56 0.6 1.3
+ 56 0.6 1.325
+ 56 0.6 1.35
+ 56 0.6 1.375
+ 56 0.6 1.4
+ 56 0.6 1.425
+ 56 0.6 1.45
+ 56 0.6 1.475
+ 56 0.6 1.5
+ 56 0.6 1.525
+ 56 0.6 1.55
+ 56 0.6 1.575
+ 56 0.6 1.6
+ 56 0.6 1.625
+ 56 0.6 1.65
+ 56 0.6 1.675
+ 56 0.6 1.7
+ 56 0.6 1.725
+ 56 0.6 1.75
+ 56 0.6 1.775
+ 56 0.6 1.8
+ 56 0.6 1.825
+ 56 0.6 1.85
+ 56 0.6 1.875
+ 56 0.6 1.9
+ 56 0.6 1.925
+ 56 0.6 1.95
+ 56 0.6 1.975
+ 56 0.6 2.0
+ 56 0.6 2.025
+ 56 0.6 2.05
+ 56 0.6 2.075
+ 56 0.6 2.1
+ 56 0.6 2.125
+ 56 0.6 2.15
+ 56 0.6 2.175
+ 56 0.6 2.2
+ 56 0.6 2.225
+ 56 0.6 2.25
+ 56 0.6 2.275
+ 56 0.6 2.3
+ 56 0.6 2.325
+ 56 0.6 2.35
+ 56 0.6 2.375
+ 56 0.6 2.4
+ 56 0.6 2.425
+ 56 0.6 2.45
+ 56 0.6 2.475
+ 56 0.6 2.5
+ 58 0.6 1.25
+ 58 0.6 1.275
+ 58 0.6 1.3
+ 58 0.6 1.325
+ 58 0.6 1.35
+ 58 0.6 1.375
+ 58 0.6 1.4
+ 58 0.6 1.425
+ 58 0.6 1.45
+ 58 0.6 1.475
+ 58 0.6 1.5
+ 58 0.6 1.525
+ 58 0.6 1.55
+ 58 0.6 1.575
+ 58 0.6 1.6
+ 58 0.6 1.625
+ 58 0.6 1.65
+ 58 0.6 1.675
+ 58 0.6 1.7
+ 58 0.6 1.725
+ 58 0.6 1.75
+ 58 0.6 1.775
+ 58 0.6 1.8
+ 58 0.6 1.825
+ 58 0.6 1.85
+ 58 0.6 1.875
+ 58 0.6 1.9
+ 58 0.6 1.925
+ 58 0.6 1.95
+ 58 0.6 1.975
+ 58 0.6 2.0
+ 58 0.6 2.025
+ 58 0.6 2.05
+ 58 0.6 2.075
+ 58 0.6 2.1
+ 58 0.6 2.125
+ 58 0.6 2.15
+ 58 0.6 2.175
+ 58 0.6 2.2
+ 58 0.6 2.225
+ 58 0.6 2.25
+ 58 0.6 2.275
+ 58 0.6 2.3
+ 58 0.6 2.325
+ 58 0.6 2.35
+ 58 0.6 2.375
+ 58 0.6 2.4
+ 58 0.6 2.425
+ 58 0.6 2.45
+ 58 0.6 2.475
+ 58 0.6 2.5
+ 60 0.6 1.25
+ 60 0.6 1.275
+ 60 0.6 1.3
+ 60 0.6 1.325
+ 60 0.6 1.35
+ 60 0.6 1.375
+ 60 0.6 1.4
+ 60 0.6 1.425
+ 60 0.6 1.45
+ 60 0.6 1.475
+ 60 0.6 1.5
+ 60 0.6 1.525
+ 60 0.6 1.55
+ 60 0.6 1.575
+ 60 0.6 1.6
+ 60 0.6 1.625
+ 60 0.6 1.65
+ 60 0.6 1.675
+ 60 0.6 1.7
+ 60 0.6 1.725
+ 60 0.6 1.75
+ 60 0.6 1.775
+ 60 0.6 1.8
+ 60 0.6 1.825
+ 60 0.6 1.85
+ 60 0.6 1.875
+ 60 0.6 1.9
+ 60 0.6 1.925
+ 60 0.6 1.95
+ 60 0.6 1.975
+ 60 0.6 2.0
+ 60 0.6 2.025
+ 60 0.6 2.05
+ 60 0.6 2.075
+ 60 0.6 2.1
+ 60 0.6 2.125
+ 60 0.6 2.15
+ 60 0.6 2.175
+ 60 0.6 2.2
+ 60 0.6 2.225
+ 60 0.6 2.25
+ 60 0.6 2.275
+ 60 0.6 2.3
+ 60 0.6 2.325
+ 60 0.6 2.35
+ 60 0.6 2.375
+ 60 0.6 2.4
+ 60 0.6 2.425
+ 60 0.6 2.45
+ 60 0.6 2.475
+ 60 0.6 2.5
+ 62 0.6 1.25
+ 62 0.6 1.275
+ 62 0.6 1.3
+ 62 0.6 1.325
+ 62 0.6 1.35
+ 62 0.6 1.375
+ 62 0.6 1.4
+ 62 0.6 1.425
+ 62 0.6 1.45
+ 62 0.6 1.475
+ 62 0.6 1.5
+ 62 0.6 1.525
+ 62 0.6 1.55
+ 62 0.6 1.575
+ 62 0.6 1.6
+ 62 0.6 1.625
+ 62 0.6 1.65
+ 62 0.6 1.675
+ 62 0.6 1.7
+ 62 0.6 1.725
+ 62 0.6 1.75
+ 62 0.6 1.775
+ 62 0.6 1.8
+ 62 0.6 1.825
+ 62 0.6 1.85
+ 62 0.6 1.875
+ 62 0.6 1.9
+ 62 0.6 1.925
+ 62 0.6 1.95
+ 62 0.6 1.975
+ 62 0.6 2.0
+ 62 0.6 2.025
+ 62 0.6 2.05
+ 62 0.6 2.075
+ 62 0.6 2.1
+ 62 0.6 2.125
+ 62 0.6 2.15
+ 62 0.6 2.175
+ 62 0.6 2.2
+ 62 0.6 2.225
+ 62 0.6 2.25
+ 62 0.6 2.275
+ 62 0.6 2.3
+ 62 0.6 2.325
+ 62 0.6 2.35
+ 62 0.6 2.375
+ 62 0.6 2.4
+ 62 0.6 2.425
+ 62 0.6 2.45
+ 62 0.6 2.475
+ 62 0.6 2.5
+ 64 0.6 1.25
+ 64 0.6 1.275
+ 64 0.6 1.3
+ 64 0.6 1.325
+ 64 0.6 1.35
+ 64 0.6 1.375
+ 64 0.6 1.4
+ 64 0.6 1.425
+ 64 0.6 1.45
+ 64 0.6 1.475
+ 64 0.6 1.5
+ 64 0.6 1.525
+ 64 0.6 1.55
+ 64 0.6 1.575
+ 64 0.6 1.6
+ 64 0.6 1.625
+ 64 0.6 1.65
+ 64 0.6 1.675
+ 64 0.6 1.7
+ 64 0.6 1.725
+ 64 0.6 1.75
+ 64 0.6 1.775
+ 64 0.6 1.8
+ 64 0.6 1.825
+ 64 0.6 1.85
+ 64 0.6 1.875
+ 64 0.6 1.9
+ 64 0.6 1.925
+ 64 0.6 1.95
+ 64 0.6 1.975
+ 64 0.6 2.0
+ 64 0.6 2.025
+ 64 0.6 2.05
+ 64 0.6 2.075
+ 64 0.6 2.1
+ 64 0.6 2.125
+ 64 0.6 2.15
+ 64 0.6 2.175
+ 64 0.6 2.2
+ 64 0.6 2.225
+ 64 0.6 2.25
+ 64 0.6 2.275
+ 64 0.6 2.3
+ 64 0.6 2.325
+ 64 0.6 2.35
+ 64 0.6 2.375
+ 64 0.6 2.4
+ 64 0.6 2.425
+ 64 0.6 2.45
+ 64 0.6 2.475
+ 64 0.6 2.5
+ 66 0.6 1.25
+ 66 0.6 1.275
+ 66 0.6 1.3
+ 66 0.6 1.325
+ 66 0.6 1.35
+ 66 0.6 1.375
+ 66 0.6 1.4
+ 66 0.6 1.425
+ 66 0.6 1.45
+ 66 0.6 1.475
+ 66 0.6 1.5
+ 66 0.6 1.525
+ 66 0.6 1.55
+ 66 0.6 1.575
+ 66 0.6 1.6
+ 66 0.6 1.625
+ 66 0.6 1.65
+ 66 0.6 1.675
+ 66 0.6 1.7
+ 66 0.6 1.725
+ 66 0.6 1.75
+ 66 0.6 1.775
+ 66 0.6 1.8
+ 66 0.6 1.825
+ 66 0.6 1.85
+ 66 0.6 1.875
+ 66 0.6 1.9
+ 66 0.6 1.925
+ 66 0.6 1.95
+ 66 0.6 1.975
+ 66 0.6 2.0
+ 66 0.6 2.025
+ 66 0.6 2.05
+ 66 0.6 2.075
+ 66 0.6 2.1
+ 66 0.6 2.125
+ 66 0.6 2.15
+ 66 0.6 2.175
+ 66 0.6 2.2
+ 66 0.6 2.225
+ 66 0.6 2.25
+ 66 0.6 2.275
+ 66 0.6 2.3
+ 66 0.6 2.325
+ 66 0.6 2.35
+ 66 0.6 2.375
+ 66 0.6 2.4
+ 66 0.6 2.425
+ 66 0.6 2.45
+ 66 0.6 2.475
+ 66 0.6 2.5
+ 68 0.6 1.25
+ 68 0.6 1.275
+ 68 0.6 1.3
+ 68 0.6 1.325
+ 68 0.6 1.35
+ 68 0.6 1.375
+ 68 0.6 1.4
+ 68 0.6 1.425
+ 68 0.6 1.45
+ 68 0.6 1.475
+ 68 0.6 1.5
+ 68 0.6 1.525
+ 68 0.6 1.55
+ 68 0.6 1.575
+ 68 0.6 1.6
+ 68 0.6 1.625
+ 68 0.6 1.65
+ 68 0.6 1.675
+ 68 0.6 1.7
+ 68 0.6 1.725
+ 68 0.6 1.75
+ 68 0.6 1.775
+ 68 0.6 1.8
+ 68 0.6 1.825
+ 68 0.6 1.85
+ 68 0.6 1.875
+ 68 0.6 1.9
+ 68 0.6 1.925
+ 68 0.6 1.95
+ 68 0.6 1.975
+ 68 0.6 2.0
+ 68 0.6 2.025
+ 68 0.6 2.05
+ 68 0.6 2.075
+ 68 0.6 2.1
+ 68 0.6 2.125
+ 68 0.6 2.15
+ 68 0.6 2.175
+ 68 0.6 2.2
+ 68 0.6 2.225
+ 68 0.6 2.25
+ 68 0.6 2.275
+ 68 0.6 2.3
+ 68 0.6 2.325
+ 68 0.6 2.35
+ 68 0.6 2.375
+ 68 0.6 2.4
+ 68 0.6 2.425
+ 68 0.6 2.45
+ 68 0.6 2.475
+ 68 0.6 2.5
+ 70 0.6 1.25
+ 70 0.6 1.275
+ 70 0.6 1.3
+ 70 0.6 1.325
+ 70 0.6 1.35
+ 70 0.6 1.375
+ 70 0.6 1.4
+ 70 0.6 1.425
+ 70 0.6 1.45
+ 70 0.6 1.475
+ 70 0.6 1.5
+ 70 0.6 1.525
+ 70 0.6 1.55
+ 70 0.6 1.575
+ 70 0.6 1.6
+ 70 0.6 1.625
+ 70 0.6 1.65
+ 70 0.6 1.675
+ 70 0.6 1.7
+ 70 0.6 1.725
+ 70 0.6 1.75
+ 70 0.6 1.775
+ 70 0.6 1.8
+ 70 0.6 1.825
+ 70 0.6 1.85
+ 70 0.6 1.875
+ 70 0.6 1.9
+ 70 0.6 1.925
+ 70 0.6 1.95
+ 70 0.6 1.975
+ 70 0.6 2.0
+ 70 0.6 2.025
+ 70 0.6 2.05
+ 70 0.6 2.075
+ 70 0.6 2.1
+ 70 0.6 2.125
+ 70 0.6 2.15
+ 70 0.6 2.175
+ 70 0.6 2.2
+ 70 0.6 2.225
+ 70 0.6 2.25
+ 70 0.6 2.275
+ 70 0.6 2.3
+ 70 0.6 2.325
+ 70 0.6 2.35
+ 70 0.6 2.375
+ 70 0.6 2.4
+ 70 0.6 2.425
+ 70 0.6 2.45
+ 70 0.6 2.475
+ 70 0.6 2.5
+ 72 0.6 1.25
+ 72 0.6 1.275
+ 72 0.6 1.3
+ 72 0.6 1.325
+ 72 0.6 1.35
+ 72 0.6 1.375
+ 72 0.6 1.4
+ 72 0.6 1.425
+ 72 0.6 1.45
+ 72 0.6 1.475
+ 72 0.6 1.5
+ 72 0.6 1.525
+ 72 0.6 1.55
+ 72 0.6 1.575
+ 72 0.6 1.6
+ 72 0.6 1.625
+ 72 0.6 1.65
+ 72 0.6 1.675
+ 72 0.6 1.7
+ 72 0.6 1.725
+ 72 0.6 1.75
+ 72 0.6 1.775
+ 72 0.6 1.8
+ 72 0.6 1.825
+ 72 0.6 1.85
+ 72 0.6 1.875
+ 72 0.6 1.9
+ 72 0.6 1.925
+ 72 0.6 1.95
+ 72 0.6 1.975
+ 72 0.6 2.0
+ 72 0.6 2.025
+ 72 0.6 2.05
+ 72 0.6 2.075
+ 72 0.6 2.1
+ 72 0.6 2.125
+ 72 0.6 2.15
+ 72 0.6 2.175
+ 72 0.6 2.2
+ 72 0.6 2.225
+ 72 0.6 2.25
+ 72 0.6 2.275
+ 72 0.6 2.3
+ 72 0.6 2.325
+ 72 0.6 2.35
+ 72 0.6 2.375
+ 72 0.6 2.4
+ 72 0.6 2.425
+ 72 0.6 2.45
+ 72 0.6 2.475
+ 72 0.6 2.5
+ 74 0.6 1.25
+ 74 0.6 1.275
+ 74 0.6 1.3
+ 74 0.6 1.325
+ 74 0.6 1.35
+ 74 0.6 1.375
+ 74 0.6 1.4
+ 74 0.6 1.425
+ 74 0.6 1.45
+ 74 0.6 1.475
+ 74 0.6 1.5
+ 74 0.6 1.525
+ 74 0.6 1.55
+ 74 0.6 1.575
+ 74 0.6 1.6
+ 74 0.6 1.625
+ 74 0.6 1.65
+ 74 0.6 1.675
+ 74 0.6 1.7
+ 74 0.6 1.725
+ 74 0.6 1.75
+ 74 0.6 1.775
+ 74 0.6 1.8
+ 74 0.6 1.825
+ 74 0.6 1.85
+ 74 0.6 1.875
+ 74 0.6 1.9
+ 74 0.6 1.925
+ 74 0.6 1.95
+ 74 0.6 1.975
+ 74 0.6 2.0
+ 74 0.6 2.025
+ 74 0.6 2.05
+ 74 0.6 2.075
+ 74 0.6 2.1
+ 74 0.6 2.125
+ 74 0.6 2.15
+ 74 0.6 2.175
+ 74 0.6 2.2
+ 74 0.6 2.225
+ 74 0.6 2.25
+ 74 0.6 2.275
+ 74 0.6 2.3
+ 74 0.6 2.325
+ 74 0.6 2.35
+ 74 0.6 2.375
+ 74 0.6 2.4
+ 74 0.6 2.425
+ 74 0.6 2.45
+ 74 0.6 2.475
+ 74 0.6 2.5
+ 76 0.6 1.25
+ 76 0.6 1.275
+ 76 0.6 1.3
+ 76 0.6 1.325
+ 76 0.6 1.35
+ 76 0.6 1.375
+ 76 0.6 1.4
+ 76 0.6 1.425
+ 76 0.6 1.45
+ 76 0.6 1.475
+ 76 0.6 1.5
+ 76 0.6 1.525
+ 76 0.6 1.55
+ 76 0.6 1.575
+ 76 0.6 1.6
+ 76 0.6 1.625
+ 76 0.6 1.65
+ 76 0.6 1.675
+ 76 0.6 1.7
+ 76 0.6 1.725
+ 76 0.6 1.75
+ 76 0.6 1.775
+ 76 0.6 1.8
+ 76 0.6 1.825
+ 76 0.6 1.85
+ 76 0.6 1.875
+ 76 0.6 1.9
+ 76 0.6 1.925
+ 76 0.6 1.95
+ 76 0.6 1.975
+ 76 0.6 2.0
+ 76 0.6 2.025
+ 76 0.6 2.05
+ 76 0.6 2.075
+ 76 0.6 2.1
+ 76 0.6 2.125
+ 76 0.6 2.15
+ 76 0.6 2.175
+ 76 0.6 2.2
+ 76 0.6 2.225
+ 76 0.6 2.25
+ 76 0.6 2.275
+ 76 0.6 2.3
+ 76 0.6 2.325
+ 76 0.6 2.35
+ 76 0.6 2.375
+ 76 0.6 2.4
+ 76 0.6 2.425
+ 76 0.6 2.45
+ 76 0.6 2.475
+ 76 0.6 2.5
+ 78 0.6 1.25
+ 78 0.6 1.275
+ 78 0.6 1.3
+ 78 0.6 1.325
+ 78 0.6 1.35
+ 78 0.6 1.375
+ 78 0.6 1.4
+ 78 0.6 1.425
+ 78 0.6 1.45
+ 78 0.6 1.475
+ 78 0.6 1.5
+ 78 0.6 1.525
+ 78 0.6 1.55
+ 78 0.6 1.575
+ 78 0.6 1.6
+ 78 0.6 1.625
+ 78 0.6 1.65
+ 78 0.6 1.675
+ 78 0.6 1.7
+ 78 0.6 1.725
+ 78 0.6 1.75
+ 78 0.6 1.775
+ 78 0.6 1.8
+ 78 0.6 1.825
+ 78 0.6 1.85
+ 78 0.6 1.875
+ 78 0.6 1.9
+ 78 0.6 1.925
+ 78 0.6 1.95
+ 78 0.6 1.975
+ 78 0.6 2.0
+ 78 0.6 2.025
+ 78 0.6 2.05
+ 78 0.6 2.075
+ 78 0.6 2.1
+ 78 0.6 2.125
+ 78 0.6 2.15
+ 78 0.6 2.175
+ 78 0.6 2.2
+ 78 0.6 2.225
+ 78 0.6 2.25
+ 78 0.6 2.275
+ 78 0.6 2.3
+ 78 0.6 2.325
+ 78 0.6 2.35
+ 78 0.6 2.375
+ 78 0.6 2.4
+ 78 0.6 2.425
+ 78 0.6 2.45
+ 78 0.6 2.475
+ 78 0.6 2.5
+ 80 0.6 1.25
+ 80 0.6 1.275
+ 80 0.6 1.3
+ 80 0.6 1.325
+ 80 0.6 1.35
+ 80 0.6 1.375
+ 80 0.6 1.4
+ 80 0.6 1.425
+ 80 0.6 1.45
+ 80 0.6 1.475
+ 80 0.6 1.5
+ 80 0.6 1.525
+ 80 0.6 1.55
+ 80 0.6 1.575
+ 80 0.6 1.6
+ 80 0.6 1.625
+ 80 0.6 1.65
+ 80 0.6 1.675
+ 80 0.6 1.7
+ 80 0.6 1.725
+ 80 0.6 1.75
+ 80 0.6 1.775
+ 80 0.6 1.8
+ 80 0.6 1.825
+ 80 0.6 1.85
+ 80 0.6 1.875
+ 80 0.6 1.9
+ 80 0.6 1.925
+ 80 0.6 1.95
+ 80 0.6 1.975
+ 80 0.6 2.0
+ 80 0.6 2.025
+ 80 0.6 2.05
+ 80 0.6 2.075
+ 80 0.6 2.1
+ 80 0.6 2.125
+ 80 0.6 2.15
+ 80 0.6 2.175
+ 80 0.6 2.2
+ 80 0.6 2.225
+ 80 0.6 2.25
+ 80 0.6 2.275
+ 80 0.6 2.3
+ 80 0.6 2.325
+ 80 0.6 2.35
+ 80 0.6 2.375
+ 80 0.6 2.4
+ 80 0.6 2.425
+ 80 0.6 2.45
+ 80 0.6 2.475
+ 80 0.6 2.5
+ 82 0.6 1.25
+ 82 0.6 1.275
+ 82 0.6 1.3
+ 82 0.6 1.325
+ 82 0.6 1.35
+ 82 0.6 1.375
+ 82 0.6 1.4
+ 82 0.6 1.425
+ 82 0.6 1.45
+ 82 0.6 1.475
+ 82 0.6 1.5
+ 82 0.6 1.525
+ 82 0.6 1.55
+ 82 0.6 1.575
+ 82 0.6 1.6
+ 82 0.6 1.625
+ 82 0.6 1.65
+ 82 0.6 1.675
+ 82 0.6 1.7
+ 82 0.6 1.725
+ 82 0.6 1.75
+ 82 0.6 1.775
+ 82 0.6 1.8
+ 82 0.6 1.825
+ 82 0.6 1.85
+ 82 0.6 1.875
+ 82 0.6 1.9
+ 82 0.6 1.925
+ 82 0.6 1.95
+ 82 0.6 1.975
+ 82 0.6 2.0
+ 82 0.6 2.025
+ 82 0.6 2.05
+ 82 0.6 2.075
+ 82 0.6 2.1
+ 82 0.6 2.125
+ 82 0.6 2.15
+ 82 0.6 2.175
+ 82 0.6 2.2
+ 82 0.6 2.225
+ 82 0.6 2.25
+ 82 0.6 2.275
+ 82 0.6 2.3
+ 82 0.6 2.325
+ 82 0.6 2.35
+ 82 0.6 2.375
+ 82 0.6 2.4
+ 82 0.6 2.425
+ 82 0.6 2.45
+ 82 0.6 2.475
+ 82 0.6 2.5
+ 84 0.6 1.25
+ 84 0.6 1.275
+ 84 0.6 1.3
+ 84 0.6 1.325
+ 84 0.6 1.35
+ 84 0.6 1.375
+ 84 0.6 1.4
+ 84 0.6 1.425
+ 84 0.6 1.45
+ 84 0.6 1.475
+ 84 0.6 1.5
+ 84 0.6 1.525
+ 84 0.6 1.55
+ 84 0.6 1.575
+ 84 0.6 1.6
+ 84 0.6 1.625
+ 84 0.6 1.65
+ 84 0.6 1.675
+ 84 0.6 1.7
+ 84 0.6 1.725
+ 84 0.6 1.75
+ 84 0.6 1.775
+ 84 0.6 1.8
+ 84 0.6 1.825
+ 84 0.6 1.85
+ 84 0.6 1.875
+ 84 0.6 1.9
+ 84 0.6 1.925
+ 84 0.6 1.95
+ 84 0.6 1.975
+ 84 0.6 2.0
+ 84 0.6 2.025
+ 84 0.6 2.05
+ 84 0.6 2.075
+ 84 0.6 2.1
+ 84 0.6 2.125
+ 84 0.6 2.15
+ 84 0.6 2.175
+ 84 0.6 2.2
+ 84 0.6 2.225
+ 84 0.6 2.25
+ 84 0.6 2.275
+ 84 0.6 2.3
+ 84 0.6 2.325
+ 84 0.6 2.35
+ 84 0.6 2.375
+ 84 0.6 2.4
+ 84 0.6 2.425
+ 84 0.6 2.45
+ 84 0.6 2.475
+ 84 0.6 2.5
+ 86 0.6 1.25
+ 86 0.6 1.275
+ 86 0.6 1.3
+ 86 0.6 1.325
+ 86 0.6 1.35
+ 86 0.6 1.375
+ 86 0.6 1.4
+ 86 0.6 1.425
+ 86 0.6 1.45
+ 86 0.6 1.475
+ 86 0.6 1.5
+ 86 0.6 1.525
+ 86 0.6 1.55
+ 86 0.6 1.575
+ 86 0.6 1.6
+ 86 0.6 1.625
+ 86 0.6 1.65
+ 86 0.6 1.675
+ 86 0.6 1.7
+ 86 0.6 1.725
+ 86 0.6 1.75
+ 86 0.6 1.775
+ 86 0.6 1.8
+ 86 0.6 1.825
+ 86 0.6 1.85
+ 86 0.6 1.875
+ 86 0.6 1.9
+ 86 0.6 1.925
+ 86 0.6 1.95
+ 86 0.6 1.975
+ 86 0.6 2.0
+ 86 0.6 2.025
+ 86 0.6 2.05
+ 86 0.6 2.075
+ 86 0.6 2.1
+ 86 0.6 2.125
+ 86 0.6 2.15
+ 86 0.6 2.175
+ 86 0.6 2.2
+ 86 0.6 2.225
+ 86 0.6 2.25
+ 86 0.6 2.275
+ 86 0.6 2.3
+ 86 0.6 2.325
+ 86 0.6 2.35
+ 86 0.6 2.375
+ 86 0.6 2.4
+ 86 0.6 2.425
+ 86 0.6 2.45
+ 86 0.6 2.475
+ 86 0.6 2.5
+ 88 0.6 1.25
+ 88 0.6 1.275
+ 88 0.6 1.3
+ 88 0.6 1.325
+ 88 0.6 1.35
+ 88 0.6 1.375
+ 88 0.6 1.4
+ 88 0.6 1.425
+ 88 0.6 1.45
+ 88 0.6 1.475
+ 88 0.6 1.5
+ 88 0.6 1.525
+ 88 0.6 1.55
+ 88 0.6 1.575
+ 88 0.6 1.6
+ 88 0.6 1.625
+ 88 0.6 1.65
+ 88 0.6 1.675
+ 88 0.6 1.7
+ 88 0.6 1.725
+ 88 0.6 1.75
+ 88 0.6 1.775
+ 88 0.6 1.8
+ 88 0.6 1.825
+ 88 0.6 1.85
+ 88 0.6 1.875
+ 88 0.6 1.9
+ 88 0.6 1.925
+ 88 0.6 1.95
+ 88 0.6 1.975
+ 88 0.6 2.0
+ 88 0.6 2.025
+ 88 0.6 2.05
+ 88 0.6 2.075
+ 88 0.6 2.1
+ 88 0.6 2.125
+ 88 0.6 2.15
+ 88 0.6 2.175
+ 88 0.6 2.2
+ 88 0.6 2.225
+ 88 0.6 2.25
+ 88 0.6 2.275
+ 88 0.6 2.3
+ 88 0.6 2.325
+ 88 0.6 2.35
+ 88 0.6 2.375
+ 88 0.6 2.4
+ 88 0.6 2.425
+ 88 0.6 2.45
+ 88 0.6 2.475
+ 88 0.6 2.5
+ 90 0.6 1.25
+ 90 0.6 1.275
+ 90 0.6 1.3
+ 90 0.6 1.325
+ 90 0.6 1.35
+ 90 0.6 1.375
+ 90 0.6 1.4
+ 90 0.6 1.425
+ 90 0.6 1.45
+ 90 0.6 1.475
+ 90 0.6 1.5
+ 90 0.6 1.525
+ 90 0.6 1.55
+ 90 0.6 1.575
+ 90 0.6 1.6
+ 90 0.6 1.625
+ 90 0.6 1.65
+ 90 0.6 1.675
+ 90 0.6 1.7
+ 90 0.6 1.725
+ 90 0.6 1.75
+ 90 0.6 1.775
+ 90 0.6 1.8
+ 90 0.6 1.825
+ 90 0.6 1.85
+ 90 0.6 1.875
+ 90 0.6 1.9
+ 90 0.6 1.925
+ 90 0.6 1.95
+ 90 0.6 1.975
+ 90 0.6 2.0
+ 90 0.6 2.025
+ 90 0.6 2.05
+ 90 0.6 2.075
+ 90 0.6 2.1
+ 90 0.6 2.125
+ 90 0.6 2.15
+ 90 0.6 2.175
+ 90 0.6 2.2
+ 90 0.6 2.225
+ 90 0.6 2.25
+ 90 0.6 2.275
+ 90 0.6 2.3
+ 90 0.6 2.325
+ 90 0.6 2.35
+ 90 0.6 2.375
+ 90 0.6 2.4
+ 90 0.6 2.425
+ 90 0.6 2.45
+ 90 0.6 2.475
+ 90 0.6 2.5
+ 92 0.6 1.25
+ 92 0.6 1.275
+ 92 0.6 1.3
+ 92 0.6 1.325
+ 92 0.6 1.35
+ 92 0.6 1.375
+ 92 0.6 1.4
+ 92 0.6 1.425
+ 92 0.6 1.45
+ 92 0.6 1.475
+ 92 0.6 1.5
+ 92 0.6 1.525
+ 92 0.6 1.55
+ 92 0.6 1.575
+ 92 0.6 1.6
+ 92 0.6 1.625
+ 92 0.6 1.65
+ 92 0.6 1.675
+ 92 0.6 1.7
+ 92 0.6 1.725
+ 92 0.6 1.75
+ 92 0.6 1.775
+ 92 0.6 1.8
+ 92 0.6 1.825
+ 92 0.6 1.85
+ 92 0.6 1.875
+ 92 0.6 1.9
+ 92 0.6 1.925
+ 92 0.6 1.95
+ 92 0.6 1.975
+ 92 0.6 2.0
+ 92 0.6 2.025
+ 92 0.6 2.05
+ 92 0.6 2.075
+ 92 0.6 2.1
+ 92 0.6 2.125
+ 92 0.6 2.15
+ 92 0.6 2.175
+ 92 0.6 2.2
+ 92 0.6 2.225
+ 92 0.6 2.25
+ 92 0.6 2.275
+ 92 0.6 2.3
+ 92 0.6 2.325
+ 92 0.6 2.35
+ 92 0.6 2.375
+ 92 0.6 2.4
+ 92 0.6 2.425
+ 92 0.6 2.45
+ 92 0.6 2.475
+ 92 0.6 2.5
+ 94 0.6 1.25
+ 94 0.6 1.275
+ 94 0.6 1.3
+ 94 0.6 1.325
+ 94 0.6 1.35
+ 94 0.6 1.375
+ 94 0.6 1.4
+ 94 0.6 1.425
+ 94 0.6 1.45
+ 94 0.6 1.475
+ 94 0.6 1.5
+ 94 0.6 1.525
+ 94 0.6 1.55
+ 94 0.6 1.575
+ 94 0.6 1.6
+ 94 0.6 1.625
+ 94 0.6 1.65
+ 94 0.6 1.675
+ 94 0.6 1.7
+ 94 0.6 1.725
+ 94 0.6 1.75
+ 94 0.6 1.775
+ 94 0.6 1.8
+ 94 0.6 1.825
+ 94 0.6 1.85
+ 94 0.6 1.875
+ 94 0.6 1.9
+ 94 0.6 1.925
+ 94 0.6 1.95
+ 94 0.6 1.975
+ 94 0.6 2.0
+ 94 0.6 2.025
+ 94 0.6 2.05
+ 94 0.6 2.075
+ 94 0.6 2.1
+ 94 0.6 2.125
+ 94 0.6 2.15
+ 94 0.6 2.175
+ 94 0.6 2.2
+ 94 0.6 2.225
+ 94 0.6 2.25
+ 94 0.6 2.275
+ 94 0.6 2.3
+ 94 0.6 2.325
+ 94 0.6 2.35
+ 94 0.6 2.375
+ 94 0.6 2.4
+ 94 0.6 2.425
+ 94 0.6 2.45
+ 94 0.6 2.475
+ 94 0.6 2.5
+ 96 0.6 1.25
+ 96 0.6 1.275
+ 96 0.6 1.3
+ 96 0.6 1.325
+ 96 0.6 1.35
+ 96 0.6 1.375
+ 96 0.6 1.4
+ 96 0.6 1.425
+ 96 0.6 1.45
+ 96 0.6 1.475
+ 96 0.6 1.5
+ 96 0.6 1.525
+ 96 0.6 1.55
+ 96 0.6 1.575
+ 96 0.6 1.6
+ 96 0.6 1.625
+ 96 0.6 1.65
+ 96 0.6 1.675
+ 96 0.6 1.7
+ 96 0.6 1.725
+ 96 0.6 1.75
+ 96 0.6 1.775
+ 96 0.6 1.8
+ 96 0.6 1.825
+ 96 0.6 1.85
+ 96 0.6 1.875
+ 96 0.6 1.9
+ 96 0.6 1.925
+ 96 0.6 1.95
+ 96 0.6 1.975
+ 96 0.6 2.0
+ 96 0.6 2.025
+ 96 0.6 2.05
+ 96 0.6 2.075
+ 96 0.6 2.1
+ 96 0.6 2.125
+ 96 0.6 2.15
+ 96 0.6 2.175
+ 96 0.6 2.2
+ 96 0.6 2.225
+ 96 0.6 2.25
+ 96 0.6 2.275
+ 96 0.6 2.3
+ 96 0.6 2.325
+ 96 0.6 2.35
+ 96 0.6 2.375
+ 96 0.6 2.4
+ 96 0.6 2.425
+ 96 0.6 2.45
+ 96 0.6 2.475
+ 96 0.6 2.5
+ 98 0.6 1.25
+ 98 0.6 1.275
+ 98 0.6 1.3
+ 98 0.6 1.325
+ 98 0.6 1.35
+ 98 0.6 1.375
+ 98 0.6 1.4
+ 98 0.6 1.425
+ 98 0.6 1.45
+ 98 0.6 1.475
+ 98 0.6 1.5
+ 98 0.6 1.525
+ 98 0.6 1.55
+ 98 0.6 1.575
+ 98 0.6 1.6
+ 98 0.6 1.625
+ 98 0.6 1.65
+ 98 0.6 1.675
+ 98 0.6 1.7
+ 98 0.6 1.725
+ 98 0.6 1.75
+ 98 0.6 1.775
+ 98 0.6 1.8
+ 98 0.6 1.825
+ 98 0.6 1.85
+ 98 0.6 1.875
+ 98 0.6 1.9
+ 98 0.6 1.925
+ 98 0.6 1.95
+ 98 0.6 1.975
+ 98 0.6 2.0
+ 98 0.6 2.025
+ 98 0.6 2.05
+ 98 0.6 2.075
+ 98 0.6 2.1
+ 98 0.6 2.125
+ 98 0.6 2.15
+ 98 0.6 2.175
+ 98 0.6 2.2
+ 98 0.6 2.225
+ 98 0.6 2.25
+ 98 0.6 2.275
+ 98 0.6 2.3
+ 98 0.6 2.325
+ 98 0.6 2.35
+ 98 0.6 2.375
+ 98 0.6 2.4
+ 98 0.6 2.425
+ 98 0.6 2.45
+ 98 0.6 2.475
+ 98 0.6 2.5
+ 100 0.6 1.25
+ 100 0.6 1.275
+ 100 0.6 1.3
+ 100 0.6 1.325
+ 100 0.6 1.35
+ 100 0.6 1.375
+ 100 0.6 1.4
+ 100 0.6 1.425
+ 100 0.6 1.45
+ 100 0.6 1.475
+ 100 0.6 1.5
+ 100 0.6 1.525
+ 100 0.6 1.55
+ 100 0.6 1.575
+ 100 0.6 1.6
+ 100 0.6 1.625
+ 100 0.6 1.65
+ 100 0.6 1.675
+ 100 0.6 1.7
+ 100 0.6 1.725
+ 100 0.6 1.75
+ 100 0.6 1.775
+ 100 0.6 1.8
+ 100 0.6 1.825
+ 100 0.6 1.85
+ 100 0.6 1.875
+ 100 0.6 1.9
+ 100 0.6 1.925
+ 100 0.6 1.95
+ 100 0.6 1.975
+ 100 0.6 2.0
+ 100 0.6 2.025
+ 100 0.6 2.05
+ 100 0.6 2.075
+ 100 0.6 2.1
+ 100 0.6 2.125
+ 100 0.6 2.15
+ 100 0.6 2.175
+ 100 0.6 2.2
+ 100 0.6 2.225
+ 100 0.6 2.25
+ 100 0.6 2.275
+ 100 0.6 2.3
+ 100 0.6 2.325
+ 100 0.6 2.35
+ 100 0.6 2.375
+ 100 0.6 2.4
+ 100 0.6 2.425
+ 100 0.6 2.45
+ 100 0.6 2.475
+ 100 0.6 2.5
+ 0 0.7 1.25
+ 0 0.7 1.275
+ 0 0.7 1.3
+ 0 0.7 1.325
+ 0 0.7 1.35
+ 0 0.7 1.375
+ 0 0.7 1.4
+ 0 0.7 1.425
+ 0 0.7 1.45
+ 0 0.7 1.475
+ 0 0.7 1.5
+ 0 0.7 1.525
+ 0 0.7 1.55
+ 0 0.7 1.575
+ 0 0.7 1.6
+ 0 0.7 1.625
+ 0 0.7 1.65
+ 0 0.7 1.675
+ 0 0.7 1.7
+ 0 0.7 1.725
+ 0 0.7 1.75
+ 0 0.7 1.775
+ 0 0.7 1.8
+ 0 0.7 1.825
+ 0 0.7 1.85
+ 0 0.7 1.875
+ 0 0.7 1.9
+ 0 0.7 1.925
+ 0 0.7 1.95
+ 0 0.7 1.975
+ 0 0.7 2.0
+ 0 0.7 2.025
+ 0 0.7 2.05
+ 0 0.7 2.075
+ 0 0.7 2.1
+ 0 0.7 2.125
+ 0 0.7 2.15
+ 0 0.7 2.175
+ 0 0.7 2.2
+ 0 0.7 2.225
+ 0 0.7 2.25
+ 0 0.7 2.275
+ 0 0.7 2.3
+ 0 0.7 2.325
+ 0 0.7 2.35
+ 0 0.7 2.375
+ 0 0.7 2.4
+ 0 0.7 2.425
+ 0 0.7 2.45
+ 0 0.7 2.475
+ 0 0.7 2.5
+ 2 0.7 1.25
+ 2 0.7 1.275
+ 2 0.7 1.3
+ 2 0.7 1.325
+ 2 0.7 1.35
+ 2 0.7 1.375
+ 2 0.7 1.4
+ 2 0.7 1.425
+ 2 0.7 1.45
+ 2 0.7 1.475
+ 2 0.7 1.5
+ 2 0.7 1.525
+ 2 0.7 1.55
+ 2 0.7 1.575
+ 2 0.7 1.6
+ 2 0.7 1.625
+ 2 0.7 1.65
+ 2 0.7 1.675
+ 2 0.7 1.7
+ 2 0.7 1.725
+ 2 0.7 1.75
+ 2 0.7 1.775
+ 2 0.7 1.8
+ 2 0.7 1.825
+ 2 0.7 1.85
+ 2 0.7 1.875
+ 2 0.7 1.9
+ 2 0.7 1.925
+ 2 0.7 1.95
+ 2 0.7 1.975
+ 2 0.7 2.0
+ 2 0.7 2.025
+ 2 0.7 2.05
+ 2 0.7 2.075
+ 2 0.7 2.1
+ 2 0.7 2.125
+ 2 0.7 2.15
+ 2 0.7 2.175
+ 2 0.7 2.2
+ 2 0.7 2.225
+ 2 0.7 2.25
+ 2 0.7 2.275
+ 2 0.7 2.3
+ 2 0.7 2.325
+ 2 0.7 2.35
+ 2 0.7 2.375
+ 2 0.7 2.4
+ 2 0.7 2.425
+ 2 0.7 2.45
+ 2 0.7 2.475
+ 2 0.7 2.5
+ 4 0.7 1.25
+ 4 0.7 1.275
+ 4 0.7 1.3
+ 4 0.7 1.325
+ 4 0.7 1.35
+ 4 0.7 1.375
+ 4 0.7 1.4
+ 4 0.7 1.425
+ 4 0.7 1.45
+ 4 0.7 1.475
+ 4 0.7 1.5
+ 4 0.7 1.525
+ 4 0.7 1.55
+ 4 0.7 1.575
+ 4 0.7 1.6
+ 4 0.7 1.625
+ 4 0.7 1.65
+ 4 0.7 1.675
+ 4 0.7 1.7
+ 4 0.7 1.725
+ 4 0.7 1.75
+ 4 0.7 1.775
+ 4 0.7 1.8
+ 4 0.7 1.825
+ 4 0.7 1.85
+ 4 0.7 1.875
+ 4 0.7 1.9
+ 4 0.7 1.925
+ 4 0.7 1.95
+ 4 0.7 1.975
+ 4 0.7 2.0
+ 4 0.7 2.025
+ 4 0.7 2.05
+ 4 0.7 2.075
+ 4 0.7 2.1
+ 4 0.7 2.125
+ 4 0.7 2.15
+ 4 0.7 2.175
+ 4 0.7 2.2
+ 4 0.7 2.225
+ 4 0.7 2.25
+ 4 0.7 2.275
+ 4 0.7 2.3
+ 4 0.7 2.325
+ 4 0.7 2.35
+ 4 0.7 2.375
+ 4 0.7 2.4
+ 4 0.7 2.425
+ 4 0.7 2.45
+ 4 0.7 2.475
+ 4 0.7 2.5
+ 6 0.7 1.25
+ 6 0.7 1.275
+ 6 0.7 1.3
+ 6 0.7 1.325
+ 6 0.7 1.35
+ 6 0.7 1.375
+ 6 0.7 1.4
+ 6 0.7 1.425
+ 6 0.7 1.45
+ 6 0.7 1.475
+ 6 0.7 1.5
+ 6 0.7 1.525
+ 6 0.7 1.55
+ 6 0.7 1.575
+ 6 0.7 1.6
+ 6 0.7 1.625
+ 6 0.7 1.65
+ 6 0.7 1.675
+ 6 0.7 1.7
+ 6 0.7 1.725
+ 6 0.7 1.75
+ 6 0.7 1.775
+ 6 0.7 1.8
+ 6 0.7 1.825
+ 6 0.7 1.85
+ 6 0.7 1.875
+ 6 0.7 1.9
+ 6 0.7 1.925
+ 6 0.7 1.95
+ 6 0.7 1.975
+ 6 0.7 2.0
+ 6 0.7 2.025
+ 6 0.7 2.05
+ 6 0.7 2.075
+ 6 0.7 2.1
+ 6 0.7 2.125
+ 6 0.7 2.15
+ 6 0.7 2.175
+ 6 0.7 2.2
+ 6 0.7 2.225
+ 6 0.7 2.25
+ 6 0.7 2.275
+ 6 0.7 2.3
+ 6 0.7 2.325
+ 6 0.7 2.35
+ 6 0.7 2.375
+ 6 0.7 2.4
+ 6 0.7 2.425
+ 6 0.7 2.45
+ 6 0.7 2.475
+ 6 0.7 2.5
+ 8 0.7 1.25
+ 8 0.7 1.275
+ 8 0.7 1.3
+ 8 0.7 1.325
+ 8 0.7 1.35
+ 8 0.7 1.375
+ 8 0.7 1.4
+ 8 0.7 1.425
+ 8 0.7 1.45
+ 8 0.7 1.475
+ 8 0.7 1.5
+ 8 0.7 1.525
+ 8 0.7 1.55
+ 8 0.7 1.575
+ 8 0.7 1.6
+ 8 0.7 1.625
+ 8 0.7 1.65
+ 8 0.7 1.675
+ 8 0.7 1.7
+ 8 0.7 1.725
+ 8 0.7 1.75
+ 8 0.7 1.775
+ 8 0.7 1.8
+ 8 0.7 1.825
+ 8 0.7 1.85
+ 8 0.7 1.875
+ 8 0.7 1.9
+ 8 0.7 1.925
+ 8 0.7 1.95
+ 8 0.7 1.975
+ 8 0.7 2.0
+ 8 0.7 2.025
+ 8 0.7 2.05
+ 8 0.7 2.075
+ 8 0.7 2.1
+ 8 0.7 2.125
+ 8 0.7 2.15
+ 8 0.7 2.175
+ 8 0.7 2.2
+ 8 0.7 2.225
+ 8 0.7 2.25
+ 8 0.7 2.275
+ 8 0.7 2.3
+ 8 0.7 2.325
+ 8 0.7 2.35
+ 8 0.7 2.375
+ 8 0.7 2.4
+ 8 0.7 2.425
+ 8 0.7 2.45
+ 8 0.7 2.475
+ 8 0.7 2.5
+ 10 0.7 1.25
+ 10 0.7 1.275
+ 10 0.7 1.3
+ 10 0.7 1.325
+ 10 0.7 1.35
+ 10 0.7 1.375
+ 10 0.7 1.4
+ 10 0.7 1.425
+ 10 0.7 1.45
+ 10 0.7 1.475
+ 10 0.7 1.5
+ 10 0.7 1.525
+ 10 0.7 1.55
+ 10 0.7 1.575
+ 10 0.7 1.6
+ 10 0.7 1.625
+ 10 0.7 1.65
+ 10 0.7 1.675
+ 10 0.7 1.7
+ 10 0.7 1.725
+ 10 0.7 1.75
+ 10 0.7 1.775
+ 10 0.7 1.8
+ 10 0.7 1.825
+ 10 0.7 1.85
+ 10 0.7 1.875
+ 10 0.7 1.9
+ 10 0.7 1.925
+ 10 0.7 1.95
+ 10 0.7 1.975
+ 10 0.7 2.0
+ 10 0.7 2.025
+ 10 0.7 2.05
+ 10 0.7 2.075
+ 10 0.7 2.1
+ 10 0.7 2.125
+ 10 0.7 2.15
+ 10 0.7 2.175
+ 10 0.7 2.2
+ 10 0.7 2.225
+ 10 0.7 2.25
+ 10 0.7 2.275
+ 10 0.7 2.3
+ 10 0.7 2.325
+ 10 0.7 2.35
+ 10 0.7 2.375
+ 10 0.7 2.4
+ 10 0.7 2.425
+ 10 0.7 2.45
+ 10 0.7 2.475
+ 10 0.7 2.5
+ 12 0.7 1.25
+ 12 0.7 1.275
+ 12 0.7 1.3
+ 12 0.7 1.325
+ 12 0.7 1.35
+ 12 0.7 1.375
+ 12 0.7 1.4
+ 12 0.7 1.425
+ 12 0.7 1.45
+ 12 0.7 1.475
+ 12 0.7 1.5
+ 12 0.7 1.525
+ 12 0.7 1.55
+ 12 0.7 1.575
+ 12 0.7 1.6
+ 12 0.7 1.625
+ 12 0.7 1.65
+ 12 0.7 1.675
+ 12 0.7 1.7
+ 12 0.7 1.725
+ 12 0.7 1.75
+ 12 0.7 1.775
+ 12 0.7 1.8
+ 12 0.7 1.825
+ 12 0.7 1.85
+ 12 0.7 1.875
+ 12 0.7 1.9
+ 12 0.7 1.925
+ 12 0.7 1.95
+ 12 0.7 1.975
+ 12 0.7 2.0
+ 12 0.7 2.025
+ 12 0.7 2.05
+ 12 0.7 2.075
+ 12 0.7 2.1
+ 12 0.7 2.125
+ 12 0.7 2.15
+ 12 0.7 2.175
+ 12 0.7 2.2
+ 12 0.7 2.225
+ 12 0.7 2.25
+ 12 0.7 2.275
+ 12 0.7 2.3
+ 12 0.7 2.325
+ 12 0.7 2.35
+ 12 0.7 2.375
+ 12 0.7 2.4
+ 12 0.7 2.425
+ 12 0.7 2.45
+ 12 0.7 2.475
+ 12 0.7 2.5
+ 14 0.7 1.25
+ 14 0.7 1.275
+ 14 0.7 1.3
+ 14 0.7 1.325
+ 14 0.7 1.35
+ 14 0.7 1.375
+ 14 0.7 1.4
+ 14 0.7 1.425
+ 14 0.7 1.45
+ 14 0.7 1.475
+ 14 0.7 1.5
+ 14 0.7 1.525
+ 14 0.7 1.55
+ 14 0.7 1.575
+ 14 0.7 1.6
+ 14 0.7 1.625
+ 14 0.7 1.65
+ 14 0.7 1.675
+ 14 0.7 1.7
+ 14 0.7 1.725
+ 14 0.7 1.75
+ 14 0.7 1.775
+ 14 0.7 1.8
+ 14 0.7 1.825
+ 14 0.7 1.85
+ 14 0.7 1.875
+ 14 0.7 1.9
+ 14 0.7 1.925
+ 14 0.7 1.95
+ 14 0.7 1.975
+ 14 0.7 2.0
+ 14 0.7 2.025
+ 14 0.7 2.05
+ 14 0.7 2.075
+ 14 0.7 2.1
+ 14 0.7 2.125
+ 14 0.7 2.15
+ 14 0.7 2.175
+ 14 0.7 2.2
+ 14 0.7 2.225
+ 14 0.7 2.25
+ 14 0.7 2.275
+ 14 0.7 2.3
+ 14 0.7 2.325
+ 14 0.7 2.35
+ 14 0.7 2.375
+ 14 0.7 2.4
+ 14 0.7 2.425
+ 14 0.7 2.45
+ 14 0.7 2.475
+ 14 0.7 2.5
+ 16 0.7 1.25
+ 16 0.7 1.275
+ 16 0.7 1.3
+ 16 0.7 1.325
+ 16 0.7 1.35
+ 16 0.7 1.375
+ 16 0.7 1.4
+ 16 0.7 1.425
+ 16 0.7 1.45
+ 16 0.7 1.475
+ 16 0.7 1.5
+ 16 0.7 1.525
+ 16 0.7 1.55
+ 16 0.7 1.575
+ 16 0.7 1.6
+ 16 0.7 1.625
+ 16 0.7 1.65
+ 16 0.7 1.675
+ 16 0.7 1.7
+ 16 0.7 1.725
+ 16 0.7 1.75
+ 16 0.7 1.775
+ 16 0.7 1.8
+ 16 0.7 1.825
+ 16 0.7 1.85
+ 16 0.7 1.875
+ 16 0.7 1.9
+ 16 0.7 1.925
+ 16 0.7 1.95
+ 16 0.7 1.975
+ 16 0.7 2.0
+ 16 0.7 2.025
+ 16 0.7 2.05
+ 16 0.7 2.075
+ 16 0.7 2.1
+ 16 0.7 2.125
+ 16 0.7 2.15
+ 16 0.7 2.175
+ 16 0.7 2.2
+ 16 0.7 2.225
+ 16 0.7 2.25
+ 16 0.7 2.275
+ 16 0.7 2.3
+ 16 0.7 2.325
+ 16 0.7 2.35
+ 16 0.7 2.375
+ 16 0.7 2.4
+ 16 0.7 2.425
+ 16 0.7 2.45
+ 16 0.7 2.475
+ 16 0.7 2.5
+ 18 0.7 1.25
+ 18 0.7 1.275
+ 18 0.7 1.3
+ 18 0.7 1.325
+ 18 0.7 1.35
+ 18 0.7 1.375
+ 18 0.7 1.4
+ 18 0.7 1.425
+ 18 0.7 1.45
+ 18 0.7 1.475
+ 18 0.7 1.5
+ 18 0.7 1.525
+ 18 0.7 1.55
+ 18 0.7 1.575
+ 18 0.7 1.6
+ 18 0.7 1.625
+ 18 0.7 1.65
+ 18 0.7 1.675
+ 18 0.7 1.7
+ 18 0.7 1.725
+ 18 0.7 1.75
+ 18 0.7 1.775
+ 18 0.7 1.8
+ 18 0.7 1.825
+ 18 0.7 1.85
+ 18 0.7 1.875
+ 18 0.7 1.9
+ 18 0.7 1.925
+ 18 0.7 1.95
+ 18 0.7 1.975
+ 18 0.7 2.0
+ 18 0.7 2.025
+ 18 0.7 2.05
+ 18 0.7 2.075
+ 18 0.7 2.1
+ 18 0.7 2.125
+ 18 0.7 2.15
+ 18 0.7 2.175
+ 18 0.7 2.2
+ 18 0.7 2.225
+ 18 0.7 2.25
+ 18 0.7 2.275
+ 18 0.7 2.3
+ 18 0.7 2.325
+ 18 0.7 2.35
+ 18 0.7 2.375
+ 18 0.7 2.4
+ 18 0.7 2.425
+ 18 0.7 2.45
+ 18 0.7 2.475
+ 18 0.7 2.5
+ 20 0.7 1.25
+ 20 0.7 1.275
+ 20 0.7 1.3
+ 20 0.7 1.325
+ 20 0.7 1.35
+ 20 0.7 1.375
+ 20 0.7 1.4
+ 20 0.7 1.425
+ 20 0.7 1.45
+ 20 0.7 1.475
+ 20 0.7 1.5
+ 20 0.7 1.525
+ 20 0.7 1.55
+ 20 0.7 1.575
+ 20 0.7 1.6
+ 20 0.7 1.625
+ 20 0.7 1.65
+ 20 0.7 1.675
+ 20 0.7 1.7
+ 20 0.7 1.725
+ 20 0.7 1.75
+ 20 0.7 1.775
+ 20 0.7 1.8
+ 20 0.7 1.825
+ 20 0.7 1.85
+ 20 0.7 1.875
+ 20 0.7 1.9
+ 20 0.7 1.925
+ 20 0.7 1.95
+ 20 0.7 1.975
+ 20 0.7 2.0
+ 20 0.7 2.025
+ 20 0.7 2.05
+ 20 0.7 2.075
+ 20 0.7 2.1
+ 20 0.7 2.125
+ 20 0.7 2.15
+ 20 0.7 2.175
+ 20 0.7 2.2
+ 20 0.7 2.225
+ 20 0.7 2.25
+ 20 0.7 2.275
+ 20 0.7 2.3
+ 20 0.7 2.325
+ 20 0.7 2.35
+ 20 0.7 2.375
+ 20 0.7 2.4
+ 20 0.7 2.425
+ 20 0.7 2.45
+ 20 0.7 2.475
+ 20 0.7 2.5
+ 22 0.7 1.25
+ 22 0.7 1.275
+ 22 0.7 1.3
+ 22 0.7 1.325
+ 22 0.7 1.35
+ 22 0.7 1.375
+ 22 0.7 1.4
+ 22 0.7 1.425
+ 22 0.7 1.45
+ 22 0.7 1.475
+ 22 0.7 1.5
+ 22 0.7 1.525
+ 22 0.7 1.55
+ 22 0.7 1.575
+ 22 0.7 1.6
+ 22 0.7 1.625
+ 22 0.7 1.65
+ 22 0.7 1.675
+ 22 0.7 1.7
+ 22 0.7 1.725
+ 22 0.7 1.75
+ 22 0.7 1.775
+ 22 0.7 1.8
+ 22 0.7 1.825
+ 22 0.7 1.85
+ 22 0.7 1.875
+ 22 0.7 1.9
+ 22 0.7 1.925
+ 22 0.7 1.95
+ 22 0.7 1.975
+ 22 0.7 2.0
+ 22 0.7 2.025
+ 22 0.7 2.05
+ 22 0.7 2.075
+ 22 0.7 2.1
+ 22 0.7 2.125
+ 22 0.7 2.15
+ 22 0.7 2.175
+ 22 0.7 2.2
+ 22 0.7 2.225
+ 22 0.7 2.25
+ 22 0.7 2.275
+ 22 0.7 2.3
+ 22 0.7 2.325
+ 22 0.7 2.35
+ 22 0.7 2.375
+ 22 0.7 2.4
+ 22 0.7 2.425
+ 22 0.7 2.45
+ 22 0.7 2.475
+ 22 0.7 2.5
+ 24 0.7 1.25
+ 24 0.7 1.275
+ 24 0.7 1.3
+ 24 0.7 1.325
+ 24 0.7 1.35
+ 24 0.7 1.375
+ 24 0.7 1.4
+ 24 0.7 1.425
+ 24 0.7 1.45
+ 24 0.7 1.475
+ 24 0.7 1.5
+ 24 0.7 1.525
+ 24 0.7 1.55
+ 24 0.7 1.575
+ 24 0.7 1.6
+ 24 0.7 1.625
+ 24 0.7 1.65
+ 24 0.7 1.675
+ 24 0.7 1.7
+ 24 0.7 1.725
+ 24 0.7 1.75
+ 24 0.7 1.775
+ 24 0.7 1.8
+ 24 0.7 1.825
+ 24 0.7 1.85
+ 24 0.7 1.875
+ 24 0.7 1.9
+ 24 0.7 1.925
+ 24 0.7 1.95
+ 24 0.7 1.975
+ 24 0.7 2.0
+ 24 0.7 2.025
+ 24 0.7 2.05
+ 24 0.7 2.075
+ 24 0.7 2.1
+ 24 0.7 2.125
+ 24 0.7 2.15
+ 24 0.7 2.175
+ 24 0.7 2.2
+ 24 0.7 2.225
+ 24 0.7 2.25
+ 24 0.7 2.275
+ 24 0.7 2.3
+ 24 0.7 2.325
+ 24 0.7 2.35
+ 24 0.7 2.375
+ 24 0.7 2.4
+ 24 0.7 2.425
+ 24 0.7 2.45
+ 24 0.7 2.475
+ 24 0.7 2.5
+ 26 0.7 1.25
+ 26 0.7 1.275
+ 26 0.7 1.3
+ 26 0.7 1.325
+ 26 0.7 1.35
+ 26 0.7 1.375
+ 26 0.7 1.4
+ 26 0.7 1.425
+ 26 0.7 1.45
+ 26 0.7 1.475
+ 26 0.7 1.5
+ 26 0.7 1.525
+ 26 0.7 1.55
+ 26 0.7 1.575
+ 26 0.7 1.6
+ 26 0.7 1.625
+ 26 0.7 1.65
+ 26 0.7 1.675
+ 26 0.7 1.7
+ 26 0.7 1.725
+ 26 0.7 1.75
+ 26 0.7 1.775
+ 26 0.7 1.8
+ 26 0.7 1.825
+ 26 0.7 1.85
+ 26 0.7 1.875
+ 26 0.7 1.9
+ 26 0.7 1.925
+ 26 0.7 1.95
+ 26 0.7 1.975
+ 26 0.7 2.0
+ 26 0.7 2.025
+ 26 0.7 2.05
+ 26 0.7 2.075
+ 26 0.7 2.1
+ 26 0.7 2.125
+ 26 0.7 2.15
+ 26 0.7 2.175
+ 26 0.7 2.2
+ 26 0.7 2.225
+ 26 0.7 2.25
+ 26 0.7 2.275
+ 26 0.7 2.3
+ 26 0.7 2.325
+ 26 0.7 2.35
+ 26 0.7 2.375
+ 26 0.7 2.4
+ 26 0.7 2.425
+ 26 0.7 2.45
+ 26 0.7 2.475
+ 26 0.7 2.5
+ 28 0.7 1.25
+ 28 0.7 1.275
+ 28 0.7 1.3
+ 28 0.7 1.325
+ 28 0.7 1.35
+ 28 0.7 1.375
+ 28 0.7 1.4
+ 28 0.7 1.425
+ 28 0.7 1.45
+ 28 0.7 1.475
+ 28 0.7 1.5
+ 28 0.7 1.525
+ 28 0.7 1.55
+ 28 0.7 1.575
+ 28 0.7 1.6
+ 28 0.7 1.625
+ 28 0.7 1.65
+ 28 0.7 1.675
+ 28 0.7 1.7
+ 28 0.7 1.725
+ 28 0.7 1.75
+ 28 0.7 1.775
+ 28 0.7 1.8
+ 28 0.7 1.825
+ 28 0.7 1.85
+ 28 0.7 1.875
+ 28 0.7 1.9
+ 28 0.7 1.925
+ 28 0.7 1.95
+ 28 0.7 1.975
+ 28 0.7 2.0
+ 28 0.7 2.025
+ 28 0.7 2.05
+ 28 0.7 2.075
+ 28 0.7 2.1
+ 28 0.7 2.125
+ 28 0.7 2.15
+ 28 0.7 2.175
+ 28 0.7 2.2
+ 28 0.7 2.225
+ 28 0.7 2.25
+ 28 0.7 2.275
+ 28 0.7 2.3
+ 28 0.7 2.325
+ 28 0.7 2.35
+ 28 0.7 2.375
+ 28 0.7 2.4
+ 28 0.7 2.425
+ 28 0.7 2.45
+ 28 0.7 2.475
+ 28 0.7 2.5
+ 30 0.7 1.25
+ 30 0.7 1.275
+ 30 0.7 1.3
+ 30 0.7 1.325
+ 30 0.7 1.35
+ 30 0.7 1.375
+ 30 0.7 1.4
+ 30 0.7 1.425
+ 30 0.7 1.45
+ 30 0.7 1.475
+ 30 0.7 1.5
+ 30 0.7 1.525
+ 30 0.7 1.55
+ 30 0.7 1.575
+ 30 0.7 1.6
+ 30 0.7 1.625
+ 30 0.7 1.65
+ 30 0.7 1.675
+ 30 0.7 1.7
+ 30 0.7 1.725
+ 30 0.7 1.75
+ 30 0.7 1.775
+ 30 0.7 1.8
+ 30 0.7 1.825
+ 30 0.7 1.85
+ 30 0.7 1.875
+ 30 0.7 1.9
+ 30 0.7 1.925
+ 30 0.7 1.95
+ 30 0.7 1.975
+ 30 0.7 2.0
+ 30 0.7 2.025
+ 30 0.7 2.05
+ 30 0.7 2.075
+ 30 0.7 2.1
+ 30 0.7 2.125
+ 30 0.7 2.15
+ 30 0.7 2.175
+ 30 0.7 2.2
+ 30 0.7 2.225
+ 30 0.7 2.25
+ 30 0.7 2.275
+ 30 0.7 2.3
+ 30 0.7 2.325
+ 30 0.7 2.35
+ 30 0.7 2.375
+ 30 0.7 2.4
+ 30 0.7 2.425
+ 30 0.7 2.45
+ 30 0.7 2.475
+ 30 0.7 2.5
+ 32 0.7 1.25
+ 32 0.7 1.275
+ 32 0.7 1.3
+ 32 0.7 1.325
+ 32 0.7 1.35
+ 32 0.7 1.375
+ 32 0.7 1.4
+ 32 0.7 1.425
+ 32 0.7 1.45
+ 32 0.7 1.475
+ 32 0.7 1.5
+ 32 0.7 1.525
+ 32 0.7 1.55
+ 32 0.7 1.575
+ 32 0.7 1.6
+ 32 0.7 1.625
+ 32 0.7 1.65
+ 32 0.7 1.675
+ 32 0.7 1.7
+ 32 0.7 1.725
+ 32 0.7 1.75
+ 32 0.7 1.775
+ 32 0.7 1.8
+ 32 0.7 1.825
+ 32 0.7 1.85
+ 32 0.7 1.875
+ 32 0.7 1.9
+ 32 0.7 1.925
+ 32 0.7 1.95
+ 32 0.7 1.975
+ 32 0.7 2.0
+ 32 0.7 2.025
+ 32 0.7 2.05
+ 32 0.7 2.075
+ 32 0.7 2.1
+ 32 0.7 2.125
+ 32 0.7 2.15
+ 32 0.7 2.175
+ 32 0.7 2.2
+ 32 0.7 2.225
+ 32 0.7 2.25
+ 32 0.7 2.275
+ 32 0.7 2.3
+ 32 0.7 2.325
+ 32 0.7 2.35
+ 32 0.7 2.375
+ 32 0.7 2.4
+ 32 0.7 2.425
+ 32 0.7 2.45
+ 32 0.7 2.475
+ 32 0.7 2.5
+ 34 0.7 1.25
+ 34 0.7 1.275
+ 34 0.7 1.3
+ 34 0.7 1.325
+ 34 0.7 1.35
+ 34 0.7 1.375
+ 34 0.7 1.4
+ 34 0.7 1.425
+ 34 0.7 1.45
+ 34 0.7 1.475
+ 34 0.7 1.5
+ 34 0.7 1.525
+ 34 0.7 1.55
+ 34 0.7 1.575
+ 34 0.7 1.6
+ 34 0.7 1.625
+ 34 0.7 1.65
+ 34 0.7 1.675
+ 34 0.7 1.7
+ 34 0.7 1.725
+ 34 0.7 1.75
+ 34 0.7 1.775
+ 34 0.7 1.8
+ 34 0.7 1.825
+ 34 0.7 1.85
+ 34 0.7 1.875
+ 34 0.7 1.9
+ 34 0.7 1.925
+ 34 0.7 1.95
+ 34 0.7 1.975
+ 34 0.7 2.0
+ 34 0.7 2.025
+ 34 0.7 2.05
+ 34 0.7 2.075
+ 34 0.7 2.1
+ 34 0.7 2.125
+ 34 0.7 2.15
+ 34 0.7 2.175
+ 34 0.7 2.2
+ 34 0.7 2.225
+ 34 0.7 2.25
+ 34 0.7 2.275
+ 34 0.7 2.3
+ 34 0.7 2.325
+ 34 0.7 2.35
+ 34 0.7 2.375
+ 34 0.7 2.4
+ 34 0.7 2.425
+ 34 0.7 2.45
+ 34 0.7 2.475
+ 34 0.7 2.5
+ 36 0.7 1.25
+ 36 0.7 1.275
+ 36 0.7 1.3
+ 36 0.7 1.325
+ 36 0.7 1.35
+ 36 0.7 1.375
+ 36 0.7 1.4
+ 36 0.7 1.425
+ 36 0.7 1.45
+ 36 0.7 1.475
+ 36 0.7 1.5
+ 36 0.7 1.525
+ 36 0.7 1.55
+ 36 0.7 1.575
+ 36 0.7 1.6
+ 36 0.7 1.625
+ 36 0.7 1.65
+ 36 0.7 1.675
+ 36 0.7 1.7
+ 36 0.7 1.725
+ 36 0.7 1.75
+ 36 0.7 1.775
+ 36 0.7 1.8
+ 36 0.7 1.825
+ 36 0.7 1.85
+ 36 0.7 1.875
+ 36 0.7 1.9
+ 36 0.7 1.925
+ 36 0.7 1.95
+ 36 0.7 1.975
+ 36 0.7 2.0
+ 36 0.7 2.025
+ 36 0.7 2.05
+ 36 0.7 2.075
+ 36 0.7 2.1
+ 36 0.7 2.125
+ 36 0.7 2.15
+ 36 0.7 2.175
+ 36 0.7 2.2
+ 36 0.7 2.225
+ 36 0.7 2.25
+ 36 0.7 2.275
+ 36 0.7 2.3
+ 36 0.7 2.325
+ 36 0.7 2.35
+ 36 0.7 2.375
+ 36 0.7 2.4
+ 36 0.7 2.425
+ 36 0.7 2.45
+ 36 0.7 2.475
+ 36 0.7 2.5
+ 38 0.7 1.25
+ 38 0.7 1.275
+ 38 0.7 1.3
+ 38 0.7 1.325
+ 38 0.7 1.35
+ 38 0.7 1.375
+ 38 0.7 1.4
+ 38 0.7 1.425
+ 38 0.7 1.45
+ 38 0.7 1.475
+ 38 0.7 1.5
+ 38 0.7 1.525
+ 38 0.7 1.55
+ 38 0.7 1.575
+ 38 0.7 1.6
+ 38 0.7 1.625
+ 38 0.7 1.65
+ 38 0.7 1.675
+ 38 0.7 1.7
+ 38 0.7 1.725
+ 38 0.7 1.75
+ 38 0.7 1.775
+ 38 0.7 1.8
+ 38 0.7 1.825
+ 38 0.7 1.85
+ 38 0.7 1.875
+ 38 0.7 1.9
+ 38 0.7 1.925
+ 38 0.7 1.95
+ 38 0.7 1.975
+ 38 0.7 2.0
+ 38 0.7 2.025
+ 38 0.7 2.05
+ 38 0.7 2.075
+ 38 0.7 2.1
+ 38 0.7 2.125
+ 38 0.7 2.15
+ 38 0.7 2.175
+ 38 0.7 2.2
+ 38 0.7 2.225
+ 38 0.7 2.25
+ 38 0.7 2.275
+ 38 0.7 2.3
+ 38 0.7 2.325
+ 38 0.7 2.35
+ 38 0.7 2.375
+ 38 0.7 2.4
+ 38 0.7 2.425
+ 38 0.7 2.45
+ 38 0.7 2.475
+ 38 0.7 2.5
+ 40 0.7 1.25
+ 40 0.7 1.275
+ 40 0.7 1.3
+ 40 0.7 1.325
+ 40 0.7 1.35
+ 40 0.7 1.375
+ 40 0.7 1.4
+ 40 0.7 1.425
+ 40 0.7 1.45
+ 40 0.7 1.475
+ 40 0.7 1.5
+ 40 0.7 1.525
+ 40 0.7 1.55
+ 40 0.7 1.575
+ 40 0.7 1.6
+ 40 0.7 1.625
+ 40 0.7 1.65
+ 40 0.7 1.675
+ 40 0.7 1.7
+ 40 0.7 1.725
+ 40 0.7 1.75
+ 40 0.7 1.775
+ 40 0.7 1.8
+ 40 0.7 1.825
+ 40 0.7 1.85
+ 40 0.7 1.875
+ 40 0.7 1.9
+ 40 0.7 1.925
+ 40 0.7 1.95
+ 40 0.7 1.975
+ 40 0.7 2.0
+ 40 0.7 2.025
+ 40 0.7 2.05
+ 40 0.7 2.075
+ 40 0.7 2.1
+ 40 0.7 2.125
+ 40 0.7 2.15
+ 40 0.7 2.175
+ 40 0.7 2.2
+ 40 0.7 2.225
+ 40 0.7 2.25
+ 40 0.7 2.275
+ 40 0.7 2.3
+ 40 0.7 2.325
+ 40 0.7 2.35
+ 40 0.7 2.375
+ 40 0.7 2.4
+ 40 0.7 2.425
+ 40 0.7 2.45
+ 40 0.7 2.475
+ 40 0.7 2.5
+ 42 0.7 1.25
+ 42 0.7 1.275
+ 42 0.7 1.3
+ 42 0.7 1.325
+ 42 0.7 1.35
+ 42 0.7 1.375
+ 42 0.7 1.4
+ 42 0.7 1.425
+ 42 0.7 1.45
+ 42 0.7 1.475
+ 42 0.7 1.5
+ 42 0.7 1.525
+ 42 0.7 1.55
+ 42 0.7 1.575
+ 42 0.7 1.6
+ 42 0.7 1.625
+ 42 0.7 1.65
+ 42 0.7 1.675
+ 42 0.7 1.7
+ 42 0.7 1.725
+ 42 0.7 1.75
+ 42 0.7 1.775
+ 42 0.7 1.8
+ 42 0.7 1.825
+ 42 0.7 1.85
+ 42 0.7 1.875
+ 42 0.7 1.9
+ 42 0.7 1.925
+ 42 0.7 1.95
+ 42 0.7 1.975
+ 42 0.7 2.0
+ 42 0.7 2.025
+ 42 0.7 2.05
+ 42 0.7 2.075
+ 42 0.7 2.1
+ 42 0.7 2.125
+ 42 0.7 2.15
+ 42 0.7 2.175
+ 42 0.7 2.2
+ 42 0.7 2.225
+ 42 0.7 2.25
+ 42 0.7 2.275
+ 42 0.7 2.3
+ 42 0.7 2.325
+ 42 0.7 2.35
+ 42 0.7 2.375
+ 42 0.7 2.4
+ 42 0.7 2.425
+ 42 0.7 2.45
+ 42 0.7 2.475
+ 42 0.7 2.5
+ 44 0.7 1.25
+ 44 0.7 1.275
+ 44 0.7 1.3
+ 44 0.7 1.325
+ 44 0.7 1.35
+ 44 0.7 1.375
+ 44 0.7 1.4
+ 44 0.7 1.425
+ 44 0.7 1.45
+ 44 0.7 1.475
+ 44 0.7 1.5
+ 44 0.7 1.525
+ 44 0.7 1.55
+ 44 0.7 1.575
+ 44 0.7 1.6
+ 44 0.7 1.625
+ 44 0.7 1.65
+ 44 0.7 1.675
+ 44 0.7 1.7
+ 44 0.7 1.725
+ 44 0.7 1.75
+ 44 0.7 1.775
+ 44 0.7 1.8
+ 44 0.7 1.825
+ 44 0.7 1.85
+ 44 0.7 1.875
+ 44 0.7 1.9
+ 44 0.7 1.925
+ 44 0.7 1.95
+ 44 0.7 1.975
+ 44 0.7 2.0
+ 44 0.7 2.025
+ 44 0.7 2.05
+ 44 0.7 2.075
+ 44 0.7 2.1
+ 44 0.7 2.125
+ 44 0.7 2.15
+ 44 0.7 2.175
+ 44 0.7 2.2
+ 44 0.7 2.225
+ 44 0.7 2.25
+ 44 0.7 2.275
+ 44 0.7 2.3
+ 44 0.7 2.325
+ 44 0.7 2.35
+ 44 0.7 2.375
+ 44 0.7 2.4
+ 44 0.7 2.425
+ 44 0.7 2.45
+ 44 0.7 2.475
+ 44 0.7 2.5
+ 46 0.7 1.25
+ 46 0.7 1.275
+ 46 0.7 1.3
+ 46 0.7 1.325
+ 46 0.7 1.35
+ 46 0.7 1.375
+ 46 0.7 1.4
+ 46 0.7 1.425
+ 46 0.7 1.45
+ 46 0.7 1.475
+ 46 0.7 1.5
+ 46 0.7 1.525
+ 46 0.7 1.55
+ 46 0.7 1.575
+ 46 0.7 1.6
+ 46 0.7 1.625
+ 46 0.7 1.65
+ 46 0.7 1.675
+ 46 0.7 1.7
+ 46 0.7 1.725
+ 46 0.7 1.75
+ 46 0.7 1.775
+ 46 0.7 1.8
+ 46 0.7 1.825
+ 46 0.7 1.85
+ 46 0.7 1.875
+ 46 0.7 1.9
+ 46 0.7 1.925
+ 46 0.7 1.95
+ 46 0.7 1.975
+ 46 0.7 2.0
+ 46 0.7 2.025
+ 46 0.7 2.05
+ 46 0.7 2.075
+ 46 0.7 2.1
+ 46 0.7 2.125
+ 46 0.7 2.15
+ 46 0.7 2.175
+ 46 0.7 2.2
+ 46 0.7 2.225
+ 46 0.7 2.25
+ 46 0.7 2.275
+ 46 0.7 2.3
+ 46 0.7 2.325
+ 46 0.7 2.35
+ 46 0.7 2.375
+ 46 0.7 2.4
+ 46 0.7 2.425
+ 46 0.7 2.45
+ 46 0.7 2.475
+ 46 0.7 2.5
+ 48 0.7 1.25
+ 48 0.7 1.275
+ 48 0.7 1.3
+ 48 0.7 1.325
+ 48 0.7 1.35
+ 48 0.7 1.375
+ 48 0.7 1.4
+ 48 0.7 1.425
+ 48 0.7 1.45
+ 48 0.7 1.475
+ 48 0.7 1.5
+ 48 0.7 1.525
+ 48 0.7 1.55
+ 48 0.7 1.575
+ 48 0.7 1.6
+ 48 0.7 1.625
+ 48 0.7 1.65
+ 48 0.7 1.675
+ 48 0.7 1.7
+ 48 0.7 1.725
+ 48 0.7 1.75
+ 48 0.7 1.775
+ 48 0.7 1.8
+ 48 0.7 1.825
+ 48 0.7 1.85
+ 48 0.7 1.875
+ 48 0.7 1.9
+ 48 0.7 1.925
+ 48 0.7 1.95
+ 48 0.7 1.975
+ 48 0.7 2.0
+ 48 0.7 2.025
+ 48 0.7 2.05
+ 48 0.7 2.075
+ 48 0.7 2.1
+ 48 0.7 2.125
+ 48 0.7 2.15
+ 48 0.7 2.175
+ 48 0.7 2.2
+ 48 0.7 2.225
+ 48 0.7 2.25
+ 48 0.7 2.275
+ 48 0.7 2.3
+ 48 0.7 2.325
+ 48 0.7 2.35
+ 48 0.7 2.375
+ 48 0.7 2.4
+ 48 0.7 2.425
+ 48 0.7 2.45
+ 48 0.7 2.475
+ 48 0.7 2.5
+ 50 0.7 1.25
+ 50 0.7 1.275
+ 50 0.7 1.3
+ 50 0.7 1.325
+ 50 0.7 1.35
+ 50 0.7 1.375
+ 50 0.7 1.4
+ 50 0.7 1.425
+ 50 0.7 1.45
+ 50 0.7 1.475
+ 50 0.7 1.5
+ 50 0.7 1.525
+ 50 0.7 1.55
+ 50 0.7 1.575
+ 50 0.7 1.6
+ 50 0.7 1.625
+ 50 0.7 1.65
+ 50 0.7 1.675
+ 50 0.7 1.7
+ 50 0.7 1.725
+ 50 0.7 1.75
+ 50 0.7 1.775
+ 50 0.7 1.8
+ 50 0.7 1.825
+ 50 0.7 1.85
+ 50 0.7 1.875
+ 50 0.7 1.9
+ 50 0.7 1.925
+ 50 0.7 1.95
+ 50 0.7 1.975
+ 50 0.7 2.0
+ 50 0.7 2.025
+ 50 0.7 2.05
+ 50 0.7 2.075
+ 50 0.7 2.1
+ 50 0.7 2.125
+ 50 0.7 2.15
+ 50 0.7 2.175
+ 50 0.7 2.2
+ 50 0.7 2.225
+ 50 0.7 2.25
+ 50 0.7 2.275
+ 50 0.7 2.3
+ 50 0.7 2.325
+ 50 0.7 2.35
+ 50 0.7 2.375
+ 50 0.7 2.4
+ 50 0.7 2.425
+ 50 0.7 2.45
+ 50 0.7 2.475
+ 50 0.7 2.5
+ 52 0.7 1.25
+ 52 0.7 1.275
+ 52 0.7 1.3
+ 52 0.7 1.325
+ 52 0.7 1.35
+ 52 0.7 1.375
+ 52 0.7 1.4
+ 52 0.7 1.425
+ 52 0.7 1.45
+ 52 0.7 1.475
+ 52 0.7 1.5
+ 52 0.7 1.525
+ 52 0.7 1.55
+ 52 0.7 1.575
+ 52 0.7 1.6
+ 52 0.7 1.625
+ 52 0.7 1.65
+ 52 0.7 1.675
+ 52 0.7 1.7
+ 52 0.7 1.725
+ 52 0.7 1.75
+ 52 0.7 1.775
+ 52 0.7 1.8
+ 52 0.7 1.825
+ 52 0.7 1.85
+ 52 0.7 1.875
+ 52 0.7 1.9
+ 52 0.7 1.925
+ 52 0.7 1.95
+ 52 0.7 1.975
+ 52 0.7 2.0
+ 52 0.7 2.025
+ 52 0.7 2.05
+ 52 0.7 2.075
+ 52 0.7 2.1
+ 52 0.7 2.125
+ 52 0.7 2.15
+ 52 0.7 2.175
+ 52 0.7 2.2
+ 52 0.7 2.225
+ 52 0.7 2.25
+ 52 0.7 2.275
+ 52 0.7 2.3
+ 52 0.7 2.325
+ 52 0.7 2.35
+ 52 0.7 2.375
+ 52 0.7 2.4
+ 52 0.7 2.425
+ 52 0.7 2.45
+ 52 0.7 2.475
+ 52 0.7 2.5
+ 54 0.7 1.25
+ 54 0.7 1.275
+ 54 0.7 1.3
+ 54 0.7 1.325
+ 54 0.7 1.35
+ 54 0.7 1.375
+ 54 0.7 1.4
+ 54 0.7 1.425
+ 54 0.7 1.45
+ 54 0.7 1.475
+ 54 0.7 1.5
+ 54 0.7 1.525
+ 54 0.7 1.55
+ 54 0.7 1.575
+ 54 0.7 1.6
+ 54 0.7 1.625
+ 54 0.7 1.65
+ 54 0.7 1.675
+ 54 0.7 1.7
+ 54 0.7 1.725
+ 54 0.7 1.75
+ 54 0.7 1.775
+ 54 0.7 1.8
+ 54 0.7 1.825
+ 54 0.7 1.85
+ 54 0.7 1.875
+ 54 0.7 1.9
+ 54 0.7 1.925
+ 54 0.7 1.95
+ 54 0.7 1.975
+ 54 0.7 2.0
+ 54 0.7 2.025
+ 54 0.7 2.05
+ 54 0.7 2.075
+ 54 0.7 2.1
+ 54 0.7 2.125
+ 54 0.7 2.15
+ 54 0.7 2.175
+ 54 0.7 2.2
+ 54 0.7 2.225
+ 54 0.7 2.25
+ 54 0.7 2.275
+ 54 0.7 2.3
+ 54 0.7 2.325
+ 54 0.7 2.35
+ 54 0.7 2.375
+ 54 0.7 2.4
+ 54 0.7 2.425
+ 54 0.7 2.45
+ 54 0.7 2.475
+ 54 0.7 2.5
+ 56 0.7 1.25
+ 56 0.7 1.275
+ 56 0.7 1.3
+ 56 0.7 1.325
+ 56 0.7 1.35
+ 56 0.7 1.375
+ 56 0.7 1.4
+ 56 0.7 1.425
+ 56 0.7 1.45
+ 56 0.7 1.475
+ 56 0.7 1.5
+ 56 0.7 1.525
+ 56 0.7 1.55
+ 56 0.7 1.575
+ 56 0.7 1.6
+ 56 0.7 1.625
+ 56 0.7 1.65
+ 56 0.7 1.675
+ 56 0.7 1.7
+ 56 0.7 1.725
+ 56 0.7 1.75
+ 56 0.7 1.775
+ 56 0.7 1.8
+ 56 0.7 1.825
+ 56 0.7 1.85
+ 56 0.7 1.875
+ 56 0.7 1.9
+ 56 0.7 1.925
+ 56 0.7 1.95
+ 56 0.7 1.975
+ 56 0.7 2.0
+ 56 0.7 2.025
+ 56 0.7 2.05
+ 56 0.7 2.075
+ 56 0.7 2.1
+ 56 0.7 2.125
+ 56 0.7 2.15
+ 56 0.7 2.175
+ 56 0.7 2.2
+ 56 0.7 2.225
+ 56 0.7 2.25
+ 56 0.7 2.275
+ 56 0.7 2.3
+ 56 0.7 2.325
+ 56 0.7 2.35
+ 56 0.7 2.375
+ 56 0.7 2.4
+ 56 0.7 2.425
+ 56 0.7 2.45
+ 56 0.7 2.475
+ 56 0.7 2.5
+ 58 0.7 1.25
+ 58 0.7 1.275
+ 58 0.7 1.3
+ 58 0.7 1.325
+ 58 0.7 1.35
+ 58 0.7 1.375
+ 58 0.7 1.4
+ 58 0.7 1.425
+ 58 0.7 1.45
+ 58 0.7 1.475
+ 58 0.7 1.5
+ 58 0.7 1.525
+ 58 0.7 1.55
+ 58 0.7 1.575
+ 58 0.7 1.6
+ 58 0.7 1.625
+ 58 0.7 1.65
+ 58 0.7 1.675
+ 58 0.7 1.7
+ 58 0.7 1.725
+ 58 0.7 1.75
+ 58 0.7 1.775
+ 58 0.7 1.8
+ 58 0.7 1.825
+ 58 0.7 1.85
+ 58 0.7 1.875
+ 58 0.7 1.9
+ 58 0.7 1.925
+ 58 0.7 1.95
+ 58 0.7 1.975
+ 58 0.7 2.0
+ 58 0.7 2.025
+ 58 0.7 2.05
+ 58 0.7 2.075
+ 58 0.7 2.1
+ 58 0.7 2.125
+ 58 0.7 2.15
+ 58 0.7 2.175
+ 58 0.7 2.2
+ 58 0.7 2.225
+ 58 0.7 2.25
+ 58 0.7 2.275
+ 58 0.7 2.3
+ 58 0.7 2.325
+ 58 0.7 2.35
+ 58 0.7 2.375
+ 58 0.7 2.4
+ 58 0.7 2.425
+ 58 0.7 2.45
+ 58 0.7 2.475
+ 58 0.7 2.5
+ 60 0.7 1.25
+ 60 0.7 1.275
+ 60 0.7 1.3
+ 60 0.7 1.325
+ 60 0.7 1.35
+ 60 0.7 1.375
+ 60 0.7 1.4
+ 60 0.7 1.425
+ 60 0.7 1.45
+ 60 0.7 1.475
+ 60 0.7 1.5
+ 60 0.7 1.525
+ 60 0.7 1.55
+ 60 0.7 1.575
+ 60 0.7 1.6
+ 60 0.7 1.625
+ 60 0.7 1.65
+ 60 0.7 1.675
+ 60 0.7 1.7
+ 60 0.7 1.725
+ 60 0.7 1.75
+ 60 0.7 1.775
+ 60 0.7 1.8
+ 60 0.7 1.825
+ 60 0.7 1.85
+ 60 0.7 1.875
+ 60 0.7 1.9
+ 60 0.7 1.925
+ 60 0.7 1.95
+ 60 0.7 1.975
+ 60 0.7 2.0
+ 60 0.7 2.025
+ 60 0.7 2.05
+ 60 0.7 2.075
+ 60 0.7 2.1
+ 60 0.7 2.125
+ 60 0.7 2.15
+ 60 0.7 2.175
+ 60 0.7 2.2
+ 60 0.7 2.225
+ 60 0.7 2.25
+ 60 0.7 2.275
+ 60 0.7 2.3
+ 60 0.7 2.325
+ 60 0.7 2.35
+ 60 0.7 2.375
+ 60 0.7 2.4
+ 60 0.7 2.425
+ 60 0.7 2.45
+ 60 0.7 2.475
+ 60 0.7 2.5
+ 62 0.7 1.25
+ 62 0.7 1.275
+ 62 0.7 1.3
+ 62 0.7 1.325
+ 62 0.7 1.35
+ 62 0.7 1.375
+ 62 0.7 1.4
+ 62 0.7 1.425
+ 62 0.7 1.45
+ 62 0.7 1.475
+ 62 0.7 1.5
+ 62 0.7 1.525
+ 62 0.7 1.55
+ 62 0.7 1.575
+ 62 0.7 1.6
+ 62 0.7 1.625
+ 62 0.7 1.65
+ 62 0.7 1.675
+ 62 0.7 1.7
+ 62 0.7 1.725
+ 62 0.7 1.75
+ 62 0.7 1.775
+ 62 0.7 1.8
+ 62 0.7 1.825
+ 62 0.7 1.85
+ 62 0.7 1.875
+ 62 0.7 1.9
+ 62 0.7 1.925
+ 62 0.7 1.95
+ 62 0.7 1.975
+ 62 0.7 2.0
+ 62 0.7 2.025
+ 62 0.7 2.05
+ 62 0.7 2.075
+ 62 0.7 2.1
+ 62 0.7 2.125
+ 62 0.7 2.15
+ 62 0.7 2.175
+ 62 0.7 2.2
+ 62 0.7 2.225
+ 62 0.7 2.25
+ 62 0.7 2.275
+ 62 0.7 2.3
+ 62 0.7 2.325
+ 62 0.7 2.35
+ 62 0.7 2.375
+ 62 0.7 2.4
+ 62 0.7 2.425
+ 62 0.7 2.45
+ 62 0.7 2.475
+ 62 0.7 2.5
+ 64 0.7 1.25
+ 64 0.7 1.275
+ 64 0.7 1.3
+ 64 0.7 1.325
+ 64 0.7 1.35
+ 64 0.7 1.375
+ 64 0.7 1.4
+ 64 0.7 1.425
+ 64 0.7 1.45
+ 64 0.7 1.475
+ 64 0.7 1.5
+ 64 0.7 1.525
+ 64 0.7 1.55
+ 64 0.7 1.575
+ 64 0.7 1.6
+ 64 0.7 1.625
+ 64 0.7 1.65
+ 64 0.7 1.675
+ 64 0.7 1.7
+ 64 0.7 1.725
+ 64 0.7 1.75
+ 64 0.7 1.775
+ 64 0.7 1.8
+ 64 0.7 1.825
+ 64 0.7 1.85
+ 64 0.7 1.875
+ 64 0.7 1.9
+ 64 0.7 1.925
+ 64 0.7 1.95
+ 64 0.7 1.975
+ 64 0.7 2.0
+ 64 0.7 2.025
+ 64 0.7 2.05
+ 64 0.7 2.075
+ 64 0.7 2.1
+ 64 0.7 2.125
+ 64 0.7 2.15
+ 64 0.7 2.175
+ 64 0.7 2.2
+ 64 0.7 2.225
+ 64 0.7 2.25
+ 64 0.7 2.275
+ 64 0.7 2.3
+ 64 0.7 2.325
+ 64 0.7 2.35
+ 64 0.7 2.375
+ 64 0.7 2.4
+ 64 0.7 2.425
+ 64 0.7 2.45
+ 64 0.7 2.475
+ 64 0.7 2.5
+ 66 0.7 1.25
+ 66 0.7 1.275
+ 66 0.7 1.3
+ 66 0.7 1.325
+ 66 0.7 1.35
+ 66 0.7 1.375
+ 66 0.7 1.4
+ 66 0.7 1.425
+ 66 0.7 1.45
+ 66 0.7 1.475
+ 66 0.7 1.5
+ 66 0.7 1.525
+ 66 0.7 1.55
+ 66 0.7 1.575
+ 66 0.7 1.6
+ 66 0.7 1.625
+ 66 0.7 1.65
+ 66 0.7 1.675
+ 66 0.7 1.7
+ 66 0.7 1.725
+ 66 0.7 1.75
+ 66 0.7 1.775
+ 66 0.7 1.8
+ 66 0.7 1.825
+ 66 0.7 1.85
+ 66 0.7 1.875
+ 66 0.7 1.9
+ 66 0.7 1.925
+ 66 0.7 1.95
+ 66 0.7 1.975
+ 66 0.7 2.0
+ 66 0.7 2.025
+ 66 0.7 2.05
+ 66 0.7 2.075
+ 66 0.7 2.1
+ 66 0.7 2.125
+ 66 0.7 2.15
+ 66 0.7 2.175
+ 66 0.7 2.2
+ 66 0.7 2.225
+ 66 0.7 2.25
+ 66 0.7 2.275
+ 66 0.7 2.3
+ 66 0.7 2.325
+ 66 0.7 2.35
+ 66 0.7 2.375
+ 66 0.7 2.4
+ 66 0.7 2.425
+ 66 0.7 2.45
+ 66 0.7 2.475
+ 66 0.7 2.5
+ 68 0.7 1.25
+ 68 0.7 1.275
+ 68 0.7 1.3
+ 68 0.7 1.325
+ 68 0.7 1.35
+ 68 0.7 1.375
+ 68 0.7 1.4
+ 68 0.7 1.425
+ 68 0.7 1.45
+ 68 0.7 1.475
+ 68 0.7 1.5
+ 68 0.7 1.525
+ 68 0.7 1.55
+ 68 0.7 1.575
+ 68 0.7 1.6
+ 68 0.7 1.625
+ 68 0.7 1.65
+ 68 0.7 1.675
+ 68 0.7 1.7
+ 68 0.7 1.725
+ 68 0.7 1.75
+ 68 0.7 1.775
+ 68 0.7 1.8
+ 68 0.7 1.825
+ 68 0.7 1.85
+ 68 0.7 1.875
+ 68 0.7 1.9
+ 68 0.7 1.925
+ 68 0.7 1.95
+ 68 0.7 1.975
+ 68 0.7 2.0
+ 68 0.7 2.025
+ 68 0.7 2.05
+ 68 0.7 2.075
+ 68 0.7 2.1
+ 68 0.7 2.125
+ 68 0.7 2.15
+ 68 0.7 2.175
+ 68 0.7 2.2
+ 68 0.7 2.225
+ 68 0.7 2.25
+ 68 0.7 2.275
+ 68 0.7 2.3
+ 68 0.7 2.325
+ 68 0.7 2.35
+ 68 0.7 2.375
+ 68 0.7 2.4
+ 68 0.7 2.425
+ 68 0.7 2.45
+ 68 0.7 2.475
+ 68 0.7 2.5
+ 70 0.7 1.25
+ 70 0.7 1.275
+ 70 0.7 1.3
+ 70 0.7 1.325
+ 70 0.7 1.35
+ 70 0.7 1.375
+ 70 0.7 1.4
+ 70 0.7 1.425
+ 70 0.7 1.45
+ 70 0.7 1.475
+ 70 0.7 1.5
+ 70 0.7 1.525
+ 70 0.7 1.55
+ 70 0.7 1.575
+ 70 0.7 1.6
+ 70 0.7 1.625
+ 70 0.7 1.65
+ 70 0.7 1.675
+ 70 0.7 1.7
+ 70 0.7 1.725
+ 70 0.7 1.75
+ 70 0.7 1.775
+ 70 0.7 1.8
+ 70 0.7 1.825
+ 70 0.7 1.85
+ 70 0.7 1.875
+ 70 0.7 1.9
+ 70 0.7 1.925
+ 70 0.7 1.95
+ 70 0.7 1.975
+ 70 0.7 2.0
+ 70 0.7 2.025
+ 70 0.7 2.05
+ 70 0.7 2.075
+ 70 0.7 2.1
+ 70 0.7 2.125
+ 70 0.7 2.15
+ 70 0.7 2.175
+ 70 0.7 2.2
+ 70 0.7 2.225
+ 70 0.7 2.25
+ 70 0.7 2.275
+ 70 0.7 2.3
+ 70 0.7 2.325
+ 70 0.7 2.35
+ 70 0.7 2.375
+ 70 0.7 2.4
+ 70 0.7 2.425
+ 70 0.7 2.45
+ 70 0.7 2.475
+ 70 0.7 2.5
+ 72 0.7 1.25
+ 72 0.7 1.275
+ 72 0.7 1.3
+ 72 0.7 1.325
+ 72 0.7 1.35
+ 72 0.7 1.375
+ 72 0.7 1.4
+ 72 0.7 1.425
+ 72 0.7 1.45
+ 72 0.7 1.475
+ 72 0.7 1.5
+ 72 0.7 1.525
+ 72 0.7 1.55
+ 72 0.7 1.575
+ 72 0.7 1.6
+ 72 0.7 1.625
+ 72 0.7 1.65
+ 72 0.7 1.675
+ 72 0.7 1.7
+ 72 0.7 1.725
+ 72 0.7 1.75
+ 72 0.7 1.775
+ 72 0.7 1.8
+ 72 0.7 1.825
+ 72 0.7 1.85
+ 72 0.7 1.875
+ 72 0.7 1.9
+ 72 0.7 1.925
+ 72 0.7 1.95
+ 72 0.7 1.975
+ 72 0.7 2.0
+ 72 0.7 2.025
+ 72 0.7 2.05
+ 72 0.7 2.075
+ 72 0.7 2.1
+ 72 0.7 2.125
+ 72 0.7 2.15
+ 72 0.7 2.175
+ 72 0.7 2.2
+ 72 0.7 2.225
+ 72 0.7 2.25
+ 72 0.7 2.275
+ 72 0.7 2.3
+ 72 0.7 2.325
+ 72 0.7 2.35
+ 72 0.7 2.375
+ 72 0.7 2.4
+ 72 0.7 2.425
+ 72 0.7 2.45
+ 72 0.7 2.475
+ 72 0.7 2.5
+ 74 0.7 1.25
+ 74 0.7 1.275
+ 74 0.7 1.3
+ 74 0.7 1.325
+ 74 0.7 1.35
+ 74 0.7 1.375
+ 74 0.7 1.4
+ 74 0.7 1.425
+ 74 0.7 1.45
+ 74 0.7 1.475
+ 74 0.7 1.5
+ 74 0.7 1.525
+ 74 0.7 1.55
+ 74 0.7 1.575
+ 74 0.7 1.6
+ 74 0.7 1.625
+ 74 0.7 1.65
+ 74 0.7 1.675
+ 74 0.7 1.7
+ 74 0.7 1.725
+ 74 0.7 1.75
+ 74 0.7 1.775
+ 74 0.7 1.8
+ 74 0.7 1.825
+ 74 0.7 1.85
+ 74 0.7 1.875
+ 74 0.7 1.9
+ 74 0.7 1.925
+ 74 0.7 1.95
+ 74 0.7 1.975
+ 74 0.7 2.0
+ 74 0.7 2.025
+ 74 0.7 2.05
+ 74 0.7 2.075
+ 74 0.7 2.1
+ 74 0.7 2.125
+ 74 0.7 2.15
+ 74 0.7 2.175
+ 74 0.7 2.2
+ 74 0.7 2.225
+ 74 0.7 2.25
+ 74 0.7 2.275
+ 74 0.7 2.3
+ 74 0.7 2.325
+ 74 0.7 2.35
+ 74 0.7 2.375
+ 74 0.7 2.4
+ 74 0.7 2.425
+ 74 0.7 2.45
+ 74 0.7 2.475
+ 74 0.7 2.5
+ 76 0.7 1.25
+ 76 0.7 1.275
+ 76 0.7 1.3
+ 76 0.7 1.325
+ 76 0.7 1.35
+ 76 0.7 1.375
+ 76 0.7 1.4
+ 76 0.7 1.425
+ 76 0.7 1.45
+ 76 0.7 1.475
+ 76 0.7 1.5
+ 76 0.7 1.525
+ 76 0.7 1.55
+ 76 0.7 1.575
+ 76 0.7 1.6
+ 76 0.7 1.625
+ 76 0.7 1.65
+ 76 0.7 1.675
+ 76 0.7 1.7
+ 76 0.7 1.725
+ 76 0.7 1.75
+ 76 0.7 1.775
+ 76 0.7 1.8
+ 76 0.7 1.825
+ 76 0.7 1.85
+ 76 0.7 1.875
+ 76 0.7 1.9
+ 76 0.7 1.925
+ 76 0.7 1.95
+ 76 0.7 1.975
+ 76 0.7 2.0
+ 76 0.7 2.025
+ 76 0.7 2.05
+ 76 0.7 2.075
+ 76 0.7 2.1
+ 76 0.7 2.125
+ 76 0.7 2.15
+ 76 0.7 2.175
+ 76 0.7 2.2
+ 76 0.7 2.225
+ 76 0.7 2.25
+ 76 0.7 2.275
+ 76 0.7 2.3
+ 76 0.7 2.325
+ 76 0.7 2.35
+ 76 0.7 2.375
+ 76 0.7 2.4
+ 76 0.7 2.425
+ 76 0.7 2.45
+ 76 0.7 2.475
+ 76 0.7 2.5
+ 78 0.7 1.25
+ 78 0.7 1.275
+ 78 0.7 1.3
+ 78 0.7 1.325
+ 78 0.7 1.35
+ 78 0.7 1.375
+ 78 0.7 1.4
+ 78 0.7 1.425
+ 78 0.7 1.45
+ 78 0.7 1.475
+ 78 0.7 1.5
+ 78 0.7 1.525
+ 78 0.7 1.55
+ 78 0.7 1.575
+ 78 0.7 1.6
+ 78 0.7 1.625
+ 78 0.7 1.65
+ 78 0.7 1.675
+ 78 0.7 1.7
+ 78 0.7 1.725
+ 78 0.7 1.75
+ 78 0.7 1.775
+ 78 0.7 1.8
+ 78 0.7 1.825
+ 78 0.7 1.85
+ 78 0.7 1.875
+ 78 0.7 1.9
+ 78 0.7 1.925
+ 78 0.7 1.95
+ 78 0.7 1.975
+ 78 0.7 2.0
+ 78 0.7 2.025
+ 78 0.7 2.05
+ 78 0.7 2.075
+ 78 0.7 2.1
+ 78 0.7 2.125
+ 78 0.7 2.15
+ 78 0.7 2.175
+ 78 0.7 2.2
+ 78 0.7 2.225
+ 78 0.7 2.25
+ 78 0.7 2.275
+ 78 0.7 2.3
+ 78 0.7 2.325
+ 78 0.7 2.35
+ 78 0.7 2.375
+ 78 0.7 2.4
+ 78 0.7 2.425
+ 78 0.7 2.45
+ 78 0.7 2.475
+ 78 0.7 2.5
+ 80 0.7 1.25
+ 80 0.7 1.275
+ 80 0.7 1.3
+ 80 0.7 1.325
+ 80 0.7 1.35
+ 80 0.7 1.375
+ 80 0.7 1.4
+ 80 0.7 1.425
+ 80 0.7 1.45
+ 80 0.7 1.475
+ 80 0.7 1.5
+ 80 0.7 1.525
+ 80 0.7 1.55
+ 80 0.7 1.575
+ 80 0.7 1.6
+ 80 0.7 1.625
+ 80 0.7 1.65
+ 80 0.7 1.675
+ 80 0.7 1.7
+ 80 0.7 1.725
+ 80 0.7 1.75
+ 80 0.7 1.775
+ 80 0.7 1.8
+ 80 0.7 1.825
+ 80 0.7 1.85
+ 80 0.7 1.875
+ 80 0.7 1.9
+ 80 0.7 1.925
+ 80 0.7 1.95
+ 80 0.7 1.975
+ 80 0.7 2.0
+ 80 0.7 2.025
+ 80 0.7 2.05
+ 80 0.7 2.075
+ 80 0.7 2.1
+ 80 0.7 2.125
+ 80 0.7 2.15
+ 80 0.7 2.175
+ 80 0.7 2.2
+ 80 0.7 2.225
+ 80 0.7 2.25
+ 80 0.7 2.275
+ 80 0.7 2.3
+ 80 0.7 2.325
+ 80 0.7 2.35
+ 80 0.7 2.375
+ 80 0.7 2.4
+ 80 0.7 2.425
+ 80 0.7 2.45
+ 80 0.7 2.475
+ 80 0.7 2.5
+ 82 0.7 1.25
+ 82 0.7 1.275
+ 82 0.7 1.3
+ 82 0.7 1.325
+ 82 0.7 1.35
+ 82 0.7 1.375
+ 82 0.7 1.4
+ 82 0.7 1.425
+ 82 0.7 1.45
+ 82 0.7 1.475
+ 82 0.7 1.5
+ 82 0.7 1.525
+ 82 0.7 1.55
+ 82 0.7 1.575
+ 82 0.7 1.6
+ 82 0.7 1.625
+ 82 0.7 1.65
+ 82 0.7 1.675
+ 82 0.7 1.7
+ 82 0.7 1.725
+ 82 0.7 1.75
+ 82 0.7 1.775
+ 82 0.7 1.8
+ 82 0.7 1.825
+ 82 0.7 1.85
+ 82 0.7 1.875
+ 82 0.7 1.9
+ 82 0.7 1.925
+ 82 0.7 1.95
+ 82 0.7 1.975
+ 82 0.7 2.0
+ 82 0.7 2.025
+ 82 0.7 2.05
+ 82 0.7 2.075
+ 82 0.7 2.1
+ 82 0.7 2.125
+ 82 0.7 2.15
+ 82 0.7 2.175
+ 82 0.7 2.2
+ 82 0.7 2.225
+ 82 0.7 2.25
+ 82 0.7 2.275
+ 82 0.7 2.3
+ 82 0.7 2.325
+ 82 0.7 2.35
+ 82 0.7 2.375
+ 82 0.7 2.4
+ 82 0.7 2.425
+ 82 0.7 2.45
+ 82 0.7 2.475
+ 82 0.7 2.5
+ 84 0.7 1.25
+ 84 0.7 1.275
+ 84 0.7 1.3
+ 84 0.7 1.325
+ 84 0.7 1.35
+ 84 0.7 1.375
+ 84 0.7 1.4
+ 84 0.7 1.425
+ 84 0.7 1.45
+ 84 0.7 1.475
+ 84 0.7 1.5
+ 84 0.7 1.525
+ 84 0.7 1.55
+ 84 0.7 1.575
+ 84 0.7 1.6
+ 84 0.7 1.625
+ 84 0.7 1.65
+ 84 0.7 1.675
+ 84 0.7 1.7
+ 84 0.7 1.725
+ 84 0.7 1.75
+ 84 0.7 1.775
+ 84 0.7 1.8
+ 84 0.7 1.825
+ 84 0.7 1.85
+ 84 0.7 1.875
+ 84 0.7 1.9
+ 84 0.7 1.925
+ 84 0.7 1.95
+ 84 0.7 1.975
+ 84 0.7 2.0
+ 84 0.7 2.025
+ 84 0.7 2.05
+ 84 0.7 2.075
+ 84 0.7 2.1
+ 84 0.7 2.125
+ 84 0.7 2.15
+ 84 0.7 2.175
+ 84 0.7 2.2
+ 84 0.7 2.225
+ 84 0.7 2.25
+ 84 0.7 2.275
+ 84 0.7 2.3
+ 84 0.7 2.325
+ 84 0.7 2.35
+ 84 0.7 2.375
+ 84 0.7 2.4
+ 84 0.7 2.425
+ 84 0.7 2.45
+ 84 0.7 2.475
+ 84 0.7 2.5
+ 86 0.7 1.25
+ 86 0.7 1.275
+ 86 0.7 1.3
+ 86 0.7 1.325
+ 86 0.7 1.35
+ 86 0.7 1.375
+ 86 0.7 1.4
+ 86 0.7 1.425
+ 86 0.7 1.45
+ 86 0.7 1.475
+ 86 0.7 1.5
+ 86 0.7 1.525
+ 86 0.7 1.55
+ 86 0.7 1.575
+ 86 0.7 1.6
+ 86 0.7 1.625
+ 86 0.7 1.65
+ 86 0.7 1.675
+ 86 0.7 1.7
+ 86 0.7 1.725
+ 86 0.7 1.75
+ 86 0.7 1.775
+ 86 0.7 1.8
+ 86 0.7 1.825
+ 86 0.7 1.85
+ 86 0.7 1.875
+ 86 0.7 1.9
+ 86 0.7 1.925
+ 86 0.7 1.95
+ 86 0.7 1.975
+ 86 0.7 2.0
+ 86 0.7 2.025
+ 86 0.7 2.05
+ 86 0.7 2.075
+ 86 0.7 2.1
+ 86 0.7 2.125
+ 86 0.7 2.15
+ 86 0.7 2.175
+ 86 0.7 2.2
+ 86 0.7 2.225
+ 86 0.7 2.25
+ 86 0.7 2.275
+ 86 0.7 2.3
+ 86 0.7 2.325
+ 86 0.7 2.35
+ 86 0.7 2.375
+ 86 0.7 2.4
+ 86 0.7 2.425
+ 86 0.7 2.45
+ 86 0.7 2.475
+ 86 0.7 2.5
+ 88 0.7 1.25
+ 88 0.7 1.275
+ 88 0.7 1.3
+ 88 0.7 1.325
+ 88 0.7 1.35
+ 88 0.7 1.375
+ 88 0.7 1.4
+ 88 0.7 1.425
+ 88 0.7 1.45
+ 88 0.7 1.475
+ 88 0.7 1.5
+ 88 0.7 1.525
+ 88 0.7 1.55
+ 88 0.7 1.575
+ 88 0.7 1.6
+ 88 0.7 1.625
+ 88 0.7 1.65
+ 88 0.7 1.675
+ 88 0.7 1.7
+ 88 0.7 1.725
+ 88 0.7 1.75
+ 88 0.7 1.775
+ 88 0.7 1.8
+ 88 0.7 1.825
+ 88 0.7 1.85
+ 88 0.7 1.875
+ 88 0.7 1.9
+ 88 0.7 1.925
+ 88 0.7 1.95
+ 88 0.7 1.975
+ 88 0.7 2.0
+ 88 0.7 2.025
+ 88 0.7 2.05
+ 88 0.7 2.075
+ 88 0.7 2.1
+ 88 0.7 2.125
+ 88 0.7 2.15
+ 88 0.7 2.175
+ 88 0.7 2.2
+ 88 0.7 2.225
+ 88 0.7 2.25
+ 88 0.7 2.275
+ 88 0.7 2.3
+ 88 0.7 2.325
+ 88 0.7 2.35
+ 88 0.7 2.375
+ 88 0.7 2.4
+ 88 0.7 2.425
+ 88 0.7 2.45
+ 88 0.7 2.475
+ 88 0.7 2.5
+ 90 0.7 1.25
+ 90 0.7 1.275
+ 90 0.7 1.3
+ 90 0.7 1.325
+ 90 0.7 1.35
+ 90 0.7 1.375
+ 90 0.7 1.4
+ 90 0.7 1.425
+ 90 0.7 1.45
+ 90 0.7 1.475
+ 90 0.7 1.5
+ 90 0.7 1.525
+ 90 0.7 1.55
+ 90 0.7 1.575
+ 90 0.7 1.6
+ 90 0.7 1.625
+ 90 0.7 1.65
+ 90 0.7 1.675
+ 90 0.7 1.7
+ 90 0.7 1.725
+ 90 0.7 1.75
+ 90 0.7 1.775
+ 90 0.7 1.8
+ 90 0.7 1.825
+ 90 0.7 1.85
+ 90 0.7 1.875
+ 90 0.7 1.9
+ 90 0.7 1.925
+ 90 0.7 1.95
+ 90 0.7 1.975
+ 90 0.7 2.0
+ 90 0.7 2.025
+ 90 0.7 2.05
+ 90 0.7 2.075
+ 90 0.7 2.1
+ 90 0.7 2.125
+ 90 0.7 2.15
+ 90 0.7 2.175
+ 90 0.7 2.2
+ 90 0.7 2.225
+ 90 0.7 2.25
+ 90 0.7 2.275
+ 90 0.7 2.3
+ 90 0.7 2.325
+ 90 0.7 2.35
+ 90 0.7 2.375
+ 90 0.7 2.4
+ 90 0.7 2.425
+ 90 0.7 2.45
+ 90 0.7 2.475
+ 90 0.7 2.5
+ 92 0.7 1.25
+ 92 0.7 1.275
+ 92 0.7 1.3
+ 92 0.7 1.325
+ 92 0.7 1.35
+ 92 0.7 1.375
+ 92 0.7 1.4
+ 92 0.7 1.425
+ 92 0.7 1.45
+ 92 0.7 1.475
+ 92 0.7 1.5
+ 92 0.7 1.525
+ 92 0.7 1.55
+ 92 0.7 1.575
+ 92 0.7 1.6
+ 92 0.7 1.625
+ 92 0.7 1.65
+ 92 0.7 1.675
+ 92 0.7 1.7
+ 92 0.7 1.725
+ 92 0.7 1.75
+ 92 0.7 1.775
+ 92 0.7 1.8
+ 92 0.7 1.825
+ 92 0.7 1.85
+ 92 0.7 1.875
+ 92 0.7 1.9
+ 92 0.7 1.925
+ 92 0.7 1.95
+ 92 0.7 1.975
+ 92 0.7 2.0
+ 92 0.7 2.025
+ 92 0.7 2.05
+ 92 0.7 2.075
+ 92 0.7 2.1
+ 92 0.7 2.125
+ 92 0.7 2.15
+ 92 0.7 2.175
+ 92 0.7 2.2
+ 92 0.7 2.225
+ 92 0.7 2.25
+ 92 0.7 2.275
+ 92 0.7 2.3
+ 92 0.7 2.325
+ 92 0.7 2.35
+ 92 0.7 2.375
+ 92 0.7 2.4
+ 92 0.7 2.425
+ 92 0.7 2.45
+ 92 0.7 2.475
+ 92 0.7 2.5
+ 94 0.7 1.25
+ 94 0.7 1.275
+ 94 0.7 1.3
+ 94 0.7 1.325
+ 94 0.7 1.35
+ 94 0.7 1.375
+ 94 0.7 1.4
+ 94 0.7 1.425
+ 94 0.7 1.45
+ 94 0.7 1.475
+ 94 0.7 1.5
+ 94 0.7 1.525
+ 94 0.7 1.55
+ 94 0.7 1.575
+ 94 0.7 1.6
+ 94 0.7 1.625
+ 94 0.7 1.65
+ 94 0.7 1.675
+ 94 0.7 1.7
+ 94 0.7 1.725
+ 94 0.7 1.75
+ 94 0.7 1.775
+ 94 0.7 1.8
+ 94 0.7 1.825
+ 94 0.7 1.85
+ 94 0.7 1.875
+ 94 0.7 1.9
+ 94 0.7 1.925
+ 94 0.7 1.95
+ 94 0.7 1.975
+ 94 0.7 2.0
+ 94 0.7 2.025
+ 94 0.7 2.05
+ 94 0.7 2.075
+ 94 0.7 2.1
+ 94 0.7 2.125
+ 94 0.7 2.15
+ 94 0.7 2.175
+ 94 0.7 2.2
+ 94 0.7 2.225
+ 94 0.7 2.25
+ 94 0.7 2.275
+ 94 0.7 2.3
+ 94 0.7 2.325
+ 94 0.7 2.35
+ 94 0.7 2.375
+ 94 0.7 2.4
+ 94 0.7 2.425
+ 94 0.7 2.45
+ 94 0.7 2.475
+ 94 0.7 2.5
+ 96 0.7 1.25
+ 96 0.7 1.275
+ 96 0.7 1.3
+ 96 0.7 1.325
+ 96 0.7 1.35
+ 96 0.7 1.375
+ 96 0.7 1.4
+ 96 0.7 1.425
+ 96 0.7 1.45
+ 96 0.7 1.475
+ 96 0.7 1.5
+ 96 0.7 1.525
+ 96 0.7 1.55
+ 96 0.7 1.575
+ 96 0.7 1.6
+ 96 0.7 1.625
+ 96 0.7 1.65
+ 96 0.7 1.675
+ 96 0.7 1.7
+ 96 0.7 1.725
+ 96 0.7 1.75
+ 96 0.7 1.775
+ 96 0.7 1.8
+ 96 0.7 1.825
+ 96 0.7 1.85
+ 96 0.7 1.875
+ 96 0.7 1.9
+ 96 0.7 1.925
+ 96 0.7 1.95
+ 96 0.7 1.975
+ 96 0.7 2.0
+ 96 0.7 2.025
+ 96 0.7 2.05
+ 96 0.7 2.075
+ 96 0.7 2.1
+ 96 0.7 2.125
+ 96 0.7 2.15
+ 96 0.7 2.175
+ 96 0.7 2.2
+ 96 0.7 2.225
+ 96 0.7 2.25
+ 96 0.7 2.275
+ 96 0.7 2.3
+ 96 0.7 2.325
+ 96 0.7 2.35
+ 96 0.7 2.375
+ 96 0.7 2.4
+ 96 0.7 2.425
+ 96 0.7 2.45
+ 96 0.7 2.475
+ 96 0.7 2.5
+ 98 0.7 1.25
+ 98 0.7 1.275
+ 98 0.7 1.3
+ 98 0.7 1.325
+ 98 0.7 1.35
+ 98 0.7 1.375
+ 98 0.7 1.4
+ 98 0.7 1.425
+ 98 0.7 1.45
+ 98 0.7 1.475
+ 98 0.7 1.5
+ 98 0.7 1.525
+ 98 0.7 1.55
+ 98 0.7 1.575
+ 98 0.7 1.6
+ 98 0.7 1.625
+ 98 0.7 1.65
+ 98 0.7 1.675
+ 98 0.7 1.7
+ 98 0.7 1.725
+ 98 0.7 1.75
+ 98 0.7 1.775
+ 98 0.7 1.8
+ 98 0.7 1.825
+ 98 0.7 1.85
+ 98 0.7 1.875
+ 98 0.7 1.9
+ 98 0.7 1.925
+ 98 0.7 1.95
+ 98 0.7 1.975
+ 98 0.7 2.0
+ 98 0.7 2.025
+ 98 0.7 2.05
+ 98 0.7 2.075
+ 98 0.7 2.1
+ 98 0.7 2.125
+ 98 0.7 2.15
+ 98 0.7 2.175
+ 98 0.7 2.2
+ 98 0.7 2.225
+ 98 0.7 2.25
+ 98 0.7 2.275
+ 98 0.7 2.3
+ 98 0.7 2.325
+ 98 0.7 2.35
+ 98 0.7 2.375
+ 98 0.7 2.4
+ 98 0.7 2.425
+ 98 0.7 2.45
+ 98 0.7 2.475
+ 98 0.7 2.5
+ 100 0.7 1.25
+ 100 0.7 1.275
+ 100 0.7 1.3
+ 100 0.7 1.325
+ 100 0.7 1.35
+ 100 0.7 1.375
+ 100 0.7 1.4
+ 100 0.7 1.425
+ 100 0.7 1.45
+ 100 0.7 1.475
+ 100 0.7 1.5
+ 100 0.7 1.525
+ 100 0.7 1.55
+ 100 0.7 1.575
+ 100 0.7 1.6
+ 100 0.7 1.625
+ 100 0.7 1.65
+ 100 0.7 1.675
+ 100 0.7 1.7
+ 100 0.7 1.725
+ 100 0.7 1.75
+ 100 0.7 1.775
+ 100 0.7 1.8
+ 100 0.7 1.825
+ 100 0.7 1.85
+ 100 0.7 1.875
+ 100 0.7 1.9
+ 100 0.7 1.925
+ 100 0.7 1.95
+ 100 0.7 1.975
+ 100 0.7 2.0
+ 100 0.7 2.025
+ 100 0.7 2.05
+ 100 0.7 2.075
+ 100 0.7 2.1
+ 100 0.7 2.125
+ 100 0.7 2.15
+ 100 0.7 2.175
+ 100 0.7 2.2
+ 100 0.7 2.225
+ 100 0.7 2.25
+ 100 0.7 2.275
+ 100 0.7 2.3
+ 100 0.7 2.325
+ 100 0.7 2.35
+ 100 0.7 2.375
+ 100 0.7 2.4
+ 100 0.7 2.425
+ 100 0.7 2.45
+ 100 0.7 2.475
+ 100 0.7 2.5
+ 0 0.8 1.25
+ 0 0.8 1.275
+ 0 0.8 1.3
+ 0 0.8 1.325
+ 0 0.8 1.35
+ 0 0.8 1.375
+ 0 0.8 1.4
+ 0 0.8 1.425
+ 0 0.8 1.45
+ 0 0.8 1.475
+ 0 0.8 1.5
+ 0 0.8 1.525
+ 0 0.8 1.55
+ 0 0.8 1.575
+ 0 0.8 1.6
+ 0 0.8 1.625
+ 0 0.8 1.65
+ 0 0.8 1.675
+ 0 0.8 1.7
+ 0 0.8 1.725
+ 0 0.8 1.75
+ 0 0.8 1.775
+ 0 0.8 1.8
+ 0 0.8 1.825
+ 0 0.8 1.85
+ 0 0.8 1.875
+ 0 0.8 1.9
+ 0 0.8 1.925
+ 0 0.8 1.95
+ 0 0.8 1.975
+ 0 0.8 2.0
+ 0 0.8 2.025
+ 0 0.8 2.05
+ 0 0.8 2.075
+ 0 0.8 2.1
+ 0 0.8 2.125
+ 0 0.8 2.15
+ 0 0.8 2.175
+ 0 0.8 2.2
+ 0 0.8 2.225
+ 0 0.8 2.25
+ 0 0.8 2.275
+ 0 0.8 2.3
+ 0 0.8 2.325
+ 0 0.8 2.35
+ 0 0.8 2.375
+ 0 0.8 2.4
+ 0 0.8 2.425
+ 0 0.8 2.45
+ 0 0.8 2.475
+ 0 0.8 2.5
+ 2 0.8 1.25
+ 2 0.8 1.275
+ 2 0.8 1.3
+ 2 0.8 1.325
+ 2 0.8 1.35
+ 2 0.8 1.375
+ 2 0.8 1.4
+ 2 0.8 1.425
+ 2 0.8 1.45
+ 2 0.8 1.475
+ 2 0.8 1.5
+ 2 0.8 1.525
+ 2 0.8 1.55
+ 2 0.8 1.575
+ 2 0.8 1.6
+ 2 0.8 1.625
+ 2 0.8 1.65
+ 2 0.8 1.675
+ 2 0.8 1.7
+ 2 0.8 1.725
+ 2 0.8 1.75
+ 2 0.8 1.775
+ 2 0.8 1.8
+ 2 0.8 1.825
+ 2 0.8 1.85
+ 2 0.8 1.875
+ 2 0.8 1.9
+ 2 0.8 1.925
+ 2 0.8 1.95
+ 2 0.8 1.975
+ 2 0.8 2.0
+ 2 0.8 2.025
+ 2 0.8 2.05
+ 2 0.8 2.075
+ 2 0.8 2.1
+ 2 0.8 2.125
+ 2 0.8 2.15
+ 2 0.8 2.175
+ 2 0.8 2.2
+ 2 0.8 2.225
+ 2 0.8 2.25
+ 2 0.8 2.275
+ 2 0.8 2.3
+ 2 0.8 2.325
+ 2 0.8 2.35
+ 2 0.8 2.375
+ 2 0.8 2.4
+ 2 0.8 2.425
+ 2 0.8 2.45
+ 2 0.8 2.475
+ 2 0.8 2.5
+ 4 0.8 1.25
+ 4 0.8 1.275
+ 4 0.8 1.3
+ 4 0.8 1.325
+ 4 0.8 1.35
+ 4 0.8 1.375
+ 4 0.8 1.4
+ 4 0.8 1.425
+ 4 0.8 1.45
+ 4 0.8 1.475
+ 4 0.8 1.5
+ 4 0.8 1.525
+ 4 0.8 1.55
+ 4 0.8 1.575
+ 4 0.8 1.6
+ 4 0.8 1.625
+ 4 0.8 1.65
+ 4 0.8 1.675
+ 4 0.8 1.7
+ 4 0.8 1.725
+ 4 0.8 1.75
+ 4 0.8 1.775
+ 4 0.8 1.8
+ 4 0.8 1.825
+ 4 0.8 1.85
+ 4 0.8 1.875
+ 4 0.8 1.9
+ 4 0.8 1.925
+ 4 0.8 1.95
+ 4 0.8 1.975
+ 4 0.8 2.0
+ 4 0.8 2.025
+ 4 0.8 2.05
+ 4 0.8 2.075
+ 4 0.8 2.1
+ 4 0.8 2.125
+ 4 0.8 2.15
+ 4 0.8 2.175
+ 4 0.8 2.2
+ 4 0.8 2.225
+ 4 0.8 2.25
+ 4 0.8 2.275
+ 4 0.8 2.3
+ 4 0.8 2.325
+ 4 0.8 2.35
+ 4 0.8 2.375
+ 4 0.8 2.4
+ 4 0.8 2.425
+ 4 0.8 2.45
+ 4 0.8 2.475
+ 4 0.8 2.5
+ 6 0.8 1.25
+ 6 0.8 1.275
+ 6 0.8 1.3
+ 6 0.8 1.325
+ 6 0.8 1.35
+ 6 0.8 1.375
+ 6 0.8 1.4
+ 6 0.8 1.425
+ 6 0.8 1.45
+ 6 0.8 1.475
+ 6 0.8 1.5
+ 6 0.8 1.525
+ 6 0.8 1.55
+ 6 0.8 1.575
+ 6 0.8 1.6
+ 6 0.8 1.625
+ 6 0.8 1.65
+ 6 0.8 1.675
+ 6 0.8 1.7
+ 6 0.8 1.725
+ 6 0.8 1.75
+ 6 0.8 1.775
+ 6 0.8 1.8
+ 6 0.8 1.825
+ 6 0.8 1.85
+ 6 0.8 1.875
+ 6 0.8 1.9
+ 6 0.8 1.925
+ 6 0.8 1.95
+ 6 0.8 1.975
+ 6 0.8 2.0
+ 6 0.8 2.025
+ 6 0.8 2.05
+ 6 0.8 2.075
+ 6 0.8 2.1
+ 6 0.8 2.125
+ 6 0.8 2.15
+ 6 0.8 2.175
+ 6 0.8 2.2
+ 6 0.8 2.225
+ 6 0.8 2.25
+ 6 0.8 2.275
+ 6 0.8 2.3
+ 6 0.8 2.325
+ 6 0.8 2.35
+ 6 0.8 2.375
+ 6 0.8 2.4
+ 6 0.8 2.425
+ 6 0.8 2.45
+ 6 0.8 2.475
+ 6 0.8 2.5
+ 8 0.8 1.25
+ 8 0.8 1.275
+ 8 0.8 1.3
+ 8 0.8 1.325
+ 8 0.8 1.35
+ 8 0.8 1.375
+ 8 0.8 1.4
+ 8 0.8 1.425
+ 8 0.8 1.45
+ 8 0.8 1.475
+ 8 0.8 1.5
+ 8 0.8 1.525
+ 8 0.8 1.55
+ 8 0.8 1.575
+ 8 0.8 1.6
+ 8 0.8 1.625
+ 8 0.8 1.65
+ 8 0.8 1.675
+ 8 0.8 1.7
+ 8 0.8 1.725
+ 8 0.8 1.75
+ 8 0.8 1.775
+ 8 0.8 1.8
+ 8 0.8 1.825
+ 8 0.8 1.85
+ 8 0.8 1.875
+ 8 0.8 1.9
+ 8 0.8 1.925
+ 8 0.8 1.95
+ 8 0.8 1.975
+ 8 0.8 2.0
+ 8 0.8 2.025
+ 8 0.8 2.05
+ 8 0.8 2.075
+ 8 0.8 2.1
+ 8 0.8 2.125
+ 8 0.8 2.15
+ 8 0.8 2.175
+ 8 0.8 2.2
+ 8 0.8 2.225
+ 8 0.8 2.25
+ 8 0.8 2.275
+ 8 0.8 2.3
+ 8 0.8 2.325
+ 8 0.8 2.35
+ 8 0.8 2.375
+ 8 0.8 2.4
+ 8 0.8 2.425
+ 8 0.8 2.45
+ 8 0.8 2.475
+ 8 0.8 2.5
+ 10 0.8 1.25
+ 10 0.8 1.275
+ 10 0.8 1.3
+ 10 0.8 1.325
+ 10 0.8 1.35
+ 10 0.8 1.375
+ 10 0.8 1.4
+ 10 0.8 1.425
+ 10 0.8 1.45
+ 10 0.8 1.475
+ 10 0.8 1.5
+ 10 0.8 1.525
+ 10 0.8 1.55
+ 10 0.8 1.575
+ 10 0.8 1.6
+ 10 0.8 1.625
+ 10 0.8 1.65
+ 10 0.8 1.675
+ 10 0.8 1.7
+ 10 0.8 1.725
+ 10 0.8 1.75
+ 10 0.8 1.775
+ 10 0.8 1.8
+ 10 0.8 1.825
+ 10 0.8 1.85
+ 10 0.8 1.875
+ 10 0.8 1.9
+ 10 0.8 1.925
+ 10 0.8 1.95
+ 10 0.8 1.975
+ 10 0.8 2.0
+ 10 0.8 2.025
+ 10 0.8 2.05
+ 10 0.8 2.075
+ 10 0.8 2.1
+ 10 0.8 2.125
+ 10 0.8 2.15
+ 10 0.8 2.175
+ 10 0.8 2.2
+ 10 0.8 2.225
+ 10 0.8 2.25
+ 10 0.8 2.275
+ 10 0.8 2.3
+ 10 0.8 2.325
+ 10 0.8 2.35
+ 10 0.8 2.375
+ 10 0.8 2.4
+ 10 0.8 2.425
+ 10 0.8 2.45
+ 10 0.8 2.475
+ 10 0.8 2.5
+ 12 0.8 1.25
+ 12 0.8 1.275
+ 12 0.8 1.3
+ 12 0.8 1.325
+ 12 0.8 1.35
+ 12 0.8 1.375
+ 12 0.8 1.4
+ 12 0.8 1.425
+ 12 0.8 1.45
+ 12 0.8 1.475
+ 12 0.8 1.5
+ 12 0.8 1.525
+ 12 0.8 1.55
+ 12 0.8 1.575
+ 12 0.8 1.6
+ 12 0.8 1.625
+ 12 0.8 1.65
+ 12 0.8 1.675
+ 12 0.8 1.7
+ 12 0.8 1.725
+ 12 0.8 1.75
+ 12 0.8 1.775
+ 12 0.8 1.8
+ 12 0.8 1.825
+ 12 0.8 1.85
+ 12 0.8 1.875
+ 12 0.8 1.9
+ 12 0.8 1.925
+ 12 0.8 1.95
+ 12 0.8 1.975
+ 12 0.8 2.0
+ 12 0.8 2.025
+ 12 0.8 2.05
+ 12 0.8 2.075
+ 12 0.8 2.1
+ 12 0.8 2.125
+ 12 0.8 2.15
+ 12 0.8 2.175
+ 12 0.8 2.2
+ 12 0.8 2.225
+ 12 0.8 2.25
+ 12 0.8 2.275
+ 12 0.8 2.3
+ 12 0.8 2.325
+ 12 0.8 2.35
+ 12 0.8 2.375
+ 12 0.8 2.4
+ 12 0.8 2.425
+ 12 0.8 2.45
+ 12 0.8 2.475
+ 12 0.8 2.5
+ 14 0.8 1.25
+ 14 0.8 1.275
+ 14 0.8 1.3
+ 14 0.8 1.325
+ 14 0.8 1.35
+ 14 0.8 1.375
+ 14 0.8 1.4
+ 14 0.8 1.425
+ 14 0.8 1.45
+ 14 0.8 1.475
+ 14 0.8 1.5
+ 14 0.8 1.525
+ 14 0.8 1.55
+ 14 0.8 1.575
+ 14 0.8 1.6
+ 14 0.8 1.625
+ 14 0.8 1.65
+ 14 0.8 1.675
+ 14 0.8 1.7
+ 14 0.8 1.725
+ 14 0.8 1.75
+ 14 0.8 1.775
+ 14 0.8 1.8
+ 14 0.8 1.825
+ 14 0.8 1.85
+ 14 0.8 1.875
+ 14 0.8 1.9
+ 14 0.8 1.925
+ 14 0.8 1.95
+ 14 0.8 1.975
+ 14 0.8 2.0
+ 14 0.8 2.025
+ 14 0.8 2.05
+ 14 0.8 2.075
+ 14 0.8 2.1
+ 14 0.8 2.125
+ 14 0.8 2.15
+ 14 0.8 2.175
+ 14 0.8 2.2
+ 14 0.8 2.225
+ 14 0.8 2.25
+ 14 0.8 2.275
+ 14 0.8 2.3
+ 14 0.8 2.325
+ 14 0.8 2.35
+ 14 0.8 2.375
+ 14 0.8 2.4
+ 14 0.8 2.425
+ 14 0.8 2.45
+ 14 0.8 2.475
+ 14 0.8 2.5
+ 16 0.8 1.25
+ 16 0.8 1.275
+ 16 0.8 1.3
+ 16 0.8 1.325
+ 16 0.8 1.35
+ 16 0.8 1.375
+ 16 0.8 1.4
+ 16 0.8 1.425
+ 16 0.8 1.45
+ 16 0.8 1.475
+ 16 0.8 1.5
+ 16 0.8 1.525
+ 16 0.8 1.55
+ 16 0.8 1.575
+ 16 0.8 1.6
+ 16 0.8 1.625
+ 16 0.8 1.65
+ 16 0.8 1.675
+ 16 0.8 1.7
+ 16 0.8 1.725
+ 16 0.8 1.75
+ 16 0.8 1.775
+ 16 0.8 1.8
+ 16 0.8 1.825
+ 16 0.8 1.85
+ 16 0.8 1.875
+ 16 0.8 1.9
+ 16 0.8 1.925
+ 16 0.8 1.95
+ 16 0.8 1.975
+ 16 0.8 2.0
+ 16 0.8 2.025
+ 16 0.8 2.05
+ 16 0.8 2.075
+ 16 0.8 2.1
+ 16 0.8 2.125
+ 16 0.8 2.15
+ 16 0.8 2.175
+ 16 0.8 2.2
+ 16 0.8 2.225
+ 16 0.8 2.25
+ 16 0.8 2.275
+ 16 0.8 2.3
+ 16 0.8 2.325
+ 16 0.8 2.35
+ 16 0.8 2.375
+ 16 0.8 2.4
+ 16 0.8 2.425
+ 16 0.8 2.45
+ 16 0.8 2.475
+ 16 0.8 2.5
+ 18 0.8 1.25
+ 18 0.8 1.275
+ 18 0.8 1.3
+ 18 0.8 1.325
+ 18 0.8 1.35
+ 18 0.8 1.375
+ 18 0.8 1.4
+ 18 0.8 1.425
+ 18 0.8 1.45
+ 18 0.8 1.475
+ 18 0.8 1.5
+ 18 0.8 1.525
+ 18 0.8 1.55
+ 18 0.8 1.575
+ 18 0.8 1.6
+ 18 0.8 1.625
+ 18 0.8 1.65
+ 18 0.8 1.675
+ 18 0.8 1.7
+ 18 0.8 1.725
+ 18 0.8 1.75
+ 18 0.8 1.775
+ 18 0.8 1.8
+ 18 0.8 1.825
+ 18 0.8 1.85
+ 18 0.8 1.875
+ 18 0.8 1.9
+ 18 0.8 1.925
+ 18 0.8 1.95
+ 18 0.8 1.975
+ 18 0.8 2.0
+ 18 0.8 2.025
+ 18 0.8 2.05
+ 18 0.8 2.075
+ 18 0.8 2.1
+ 18 0.8 2.125
+ 18 0.8 2.15
+ 18 0.8 2.175
+ 18 0.8 2.2
+ 18 0.8 2.225
+ 18 0.8 2.25
+ 18 0.8 2.275
+ 18 0.8 2.3
+ 18 0.8 2.325
+ 18 0.8 2.35
+ 18 0.8 2.375
+ 18 0.8 2.4
+ 18 0.8 2.425
+ 18 0.8 2.45
+ 18 0.8 2.475
+ 18 0.8 2.5
+ 20 0.8 1.25
+ 20 0.8 1.275
+ 20 0.8 1.3
+ 20 0.8 1.325
+ 20 0.8 1.35
+ 20 0.8 1.375
+ 20 0.8 1.4
+ 20 0.8 1.425
+ 20 0.8 1.45
+ 20 0.8 1.475
+ 20 0.8 1.5
+ 20 0.8 1.525
+ 20 0.8 1.55
+ 20 0.8 1.575
+ 20 0.8 1.6
+ 20 0.8 1.625
+ 20 0.8 1.65
+ 20 0.8 1.675
+ 20 0.8 1.7
+ 20 0.8 1.725
+ 20 0.8 1.75
+ 20 0.8 1.775
+ 20 0.8 1.8
+ 20 0.8 1.825
+ 20 0.8 1.85
+ 20 0.8 1.875
+ 20 0.8 1.9
+ 20 0.8 1.925
+ 20 0.8 1.95
+ 20 0.8 1.975
+ 20 0.8 2.0
+ 20 0.8 2.025
+ 20 0.8 2.05
+ 20 0.8 2.075
+ 20 0.8 2.1
+ 20 0.8 2.125
+ 20 0.8 2.15
+ 20 0.8 2.175
+ 20 0.8 2.2
+ 20 0.8 2.225
+ 20 0.8 2.25
+ 20 0.8 2.275
+ 20 0.8 2.3
+ 20 0.8 2.325
+ 20 0.8 2.35
+ 20 0.8 2.375
+ 20 0.8 2.4
+ 20 0.8 2.425
+ 20 0.8 2.45
+ 20 0.8 2.475
+ 20 0.8 2.5
+ 22 0.8 1.25
+ 22 0.8 1.275
+ 22 0.8 1.3
+ 22 0.8 1.325
+ 22 0.8 1.35
+ 22 0.8 1.375
+ 22 0.8 1.4
+ 22 0.8 1.425
+ 22 0.8 1.45
+ 22 0.8 1.475
+ 22 0.8 1.5
+ 22 0.8 1.525
+ 22 0.8 1.55
+ 22 0.8 1.575
+ 22 0.8 1.6
+ 22 0.8 1.625
+ 22 0.8 1.65
+ 22 0.8 1.675
+ 22 0.8 1.7
+ 22 0.8 1.725
+ 22 0.8 1.75
+ 22 0.8 1.775
+ 22 0.8 1.8
+ 22 0.8 1.825
+ 22 0.8 1.85
+ 22 0.8 1.875
+ 22 0.8 1.9
+ 22 0.8 1.925
+ 22 0.8 1.95
+ 22 0.8 1.975
+ 22 0.8 2.0
+ 22 0.8 2.025
+ 22 0.8 2.05
+ 22 0.8 2.075
+ 22 0.8 2.1
+ 22 0.8 2.125
+ 22 0.8 2.15
+ 22 0.8 2.175
+ 22 0.8 2.2
+ 22 0.8 2.225
+ 22 0.8 2.25
+ 22 0.8 2.275
+ 22 0.8 2.3
+ 22 0.8 2.325
+ 22 0.8 2.35
+ 22 0.8 2.375
+ 22 0.8 2.4
+ 22 0.8 2.425
+ 22 0.8 2.45
+ 22 0.8 2.475
+ 22 0.8 2.5
+ 24 0.8 1.25
+ 24 0.8 1.275
+ 24 0.8 1.3
+ 24 0.8 1.325
+ 24 0.8 1.35
+ 24 0.8 1.375
+ 24 0.8 1.4
+ 24 0.8 1.425
+ 24 0.8 1.45
+ 24 0.8 1.475
+ 24 0.8 1.5
+ 24 0.8 1.525
+ 24 0.8 1.55
+ 24 0.8 1.575
+ 24 0.8 1.6
+ 24 0.8 1.625
+ 24 0.8 1.65
+ 24 0.8 1.675
+ 24 0.8 1.7
+ 24 0.8 1.725
+ 24 0.8 1.75
+ 24 0.8 1.775
+ 24 0.8 1.8
+ 24 0.8 1.825
+ 24 0.8 1.85
+ 24 0.8 1.875
+ 24 0.8 1.9
+ 24 0.8 1.925
+ 24 0.8 1.95
+ 24 0.8 1.975
+ 24 0.8 2.0
+ 24 0.8 2.025
+ 24 0.8 2.05
+ 24 0.8 2.075
+ 24 0.8 2.1
+ 24 0.8 2.125
+ 24 0.8 2.15
+ 24 0.8 2.175
+ 24 0.8 2.2
+ 24 0.8 2.225
+ 24 0.8 2.25
+ 24 0.8 2.275
+ 24 0.8 2.3
+ 24 0.8 2.325
+ 24 0.8 2.35
+ 24 0.8 2.375
+ 24 0.8 2.4
+ 24 0.8 2.425
+ 24 0.8 2.45
+ 24 0.8 2.475
+ 24 0.8 2.5
+ 26 0.8 1.25
+ 26 0.8 1.275
+ 26 0.8 1.3
+ 26 0.8 1.325
+ 26 0.8 1.35
+ 26 0.8 1.375
+ 26 0.8 1.4
+ 26 0.8 1.425
+ 26 0.8 1.45
+ 26 0.8 1.475
+ 26 0.8 1.5
+ 26 0.8 1.525
+ 26 0.8 1.55
+ 26 0.8 1.575
+ 26 0.8 1.6
+ 26 0.8 1.625
+ 26 0.8 1.65
+ 26 0.8 1.675
+ 26 0.8 1.7
+ 26 0.8 1.725
+ 26 0.8 1.75
+ 26 0.8 1.775
+ 26 0.8 1.8
+ 26 0.8 1.825
+ 26 0.8 1.85
+ 26 0.8 1.875
+ 26 0.8 1.9
+ 26 0.8 1.925
+ 26 0.8 1.95
+ 26 0.8 1.975
+ 26 0.8 2.0
+ 26 0.8 2.025
+ 26 0.8 2.05
+ 26 0.8 2.075
+ 26 0.8 2.1
+ 26 0.8 2.125
+ 26 0.8 2.15
+ 26 0.8 2.175
+ 26 0.8 2.2
+ 26 0.8 2.225
+ 26 0.8 2.25
+ 26 0.8 2.275
+ 26 0.8 2.3
+ 26 0.8 2.325
+ 26 0.8 2.35
+ 26 0.8 2.375
+ 26 0.8 2.4
+ 26 0.8 2.425
+ 26 0.8 2.45
+ 26 0.8 2.475
+ 26 0.8 2.5
+ 28 0.8 1.25
+ 28 0.8 1.275
+ 28 0.8 1.3
+ 28 0.8 1.325
+ 28 0.8 1.35
+ 28 0.8 1.375
+ 28 0.8 1.4
+ 28 0.8 1.425
+ 28 0.8 1.45
+ 28 0.8 1.475
+ 28 0.8 1.5
+ 28 0.8 1.525
+ 28 0.8 1.55
+ 28 0.8 1.575
+ 28 0.8 1.6
+ 28 0.8 1.625
+ 28 0.8 1.65
+ 28 0.8 1.675
+ 28 0.8 1.7
+ 28 0.8 1.725
+ 28 0.8 1.75
+ 28 0.8 1.775
+ 28 0.8 1.8
+ 28 0.8 1.825
+ 28 0.8 1.85
+ 28 0.8 1.875
+ 28 0.8 1.9
+ 28 0.8 1.925
+ 28 0.8 1.95
+ 28 0.8 1.975
+ 28 0.8 2.0
+ 28 0.8 2.025
+ 28 0.8 2.05
+ 28 0.8 2.075
+ 28 0.8 2.1
+ 28 0.8 2.125
+ 28 0.8 2.15
+ 28 0.8 2.175
+ 28 0.8 2.2
+ 28 0.8 2.225
+ 28 0.8 2.25
+ 28 0.8 2.275
+ 28 0.8 2.3
+ 28 0.8 2.325
+ 28 0.8 2.35
+ 28 0.8 2.375
+ 28 0.8 2.4
+ 28 0.8 2.425
+ 28 0.8 2.45
+ 28 0.8 2.475
+ 28 0.8 2.5
+ 30 0.8 1.25
+ 30 0.8 1.275
+ 30 0.8 1.3
+ 30 0.8 1.325
+ 30 0.8 1.35
+ 30 0.8 1.375
+ 30 0.8 1.4
+ 30 0.8 1.425
+ 30 0.8 1.45
+ 30 0.8 1.475
+ 30 0.8 1.5
+ 30 0.8 1.525
+ 30 0.8 1.55
+ 30 0.8 1.575
+ 30 0.8 1.6
+ 30 0.8 1.625
+ 30 0.8 1.65
+ 30 0.8 1.675
+ 30 0.8 1.7
+ 30 0.8 1.725
+ 30 0.8 1.75
+ 30 0.8 1.775
+ 30 0.8 1.8
+ 30 0.8 1.825
+ 30 0.8 1.85
+ 30 0.8 1.875
+ 30 0.8 1.9
+ 30 0.8 1.925
+ 30 0.8 1.95
+ 30 0.8 1.975
+ 30 0.8 2.0
+ 30 0.8 2.025
+ 30 0.8 2.05
+ 30 0.8 2.075
+ 30 0.8 2.1
+ 30 0.8 2.125
+ 30 0.8 2.15
+ 30 0.8 2.175
+ 30 0.8 2.2
+ 30 0.8 2.225
+ 30 0.8 2.25
+ 30 0.8 2.275
+ 30 0.8 2.3
+ 30 0.8 2.325
+ 30 0.8 2.35
+ 30 0.8 2.375
+ 30 0.8 2.4
+ 30 0.8 2.425
+ 30 0.8 2.45
+ 30 0.8 2.475
+ 30 0.8 2.5
+ 32 0.8 1.25
+ 32 0.8 1.275
+ 32 0.8 1.3
+ 32 0.8 1.325
+ 32 0.8 1.35
+ 32 0.8 1.375
+ 32 0.8 1.4
+ 32 0.8 1.425
+ 32 0.8 1.45
+ 32 0.8 1.475
+ 32 0.8 1.5
+ 32 0.8 1.525
+ 32 0.8 1.55
+ 32 0.8 1.575
+ 32 0.8 1.6
+ 32 0.8 1.625
+ 32 0.8 1.65
+ 32 0.8 1.675
+ 32 0.8 1.7
+ 32 0.8 1.725
+ 32 0.8 1.75
+ 32 0.8 1.775
+ 32 0.8 1.8
+ 32 0.8 1.825
+ 32 0.8 1.85
+ 32 0.8 1.875
+ 32 0.8 1.9
+ 32 0.8 1.925
+ 32 0.8 1.95
+ 32 0.8 1.975
+ 32 0.8 2.0
+ 32 0.8 2.025
+ 32 0.8 2.05
+ 32 0.8 2.075
+ 32 0.8 2.1
+ 32 0.8 2.125
+ 32 0.8 2.15
+ 32 0.8 2.175
+ 32 0.8 2.2
+ 32 0.8 2.225
+ 32 0.8 2.25
+ 32 0.8 2.275
+ 32 0.8 2.3
+ 32 0.8 2.325
+ 32 0.8 2.35
+ 32 0.8 2.375
+ 32 0.8 2.4
+ 32 0.8 2.425
+ 32 0.8 2.45
+ 32 0.8 2.475
+ 32 0.8 2.5
+ 34 0.8 1.25
+ 34 0.8 1.275
+ 34 0.8 1.3
+ 34 0.8 1.325
+ 34 0.8 1.35
+ 34 0.8 1.375
+ 34 0.8 1.4
+ 34 0.8 1.425
+ 34 0.8 1.45
+ 34 0.8 1.475
+ 34 0.8 1.5
+ 34 0.8 1.525
+ 34 0.8 1.55
+ 34 0.8 1.575
+ 34 0.8 1.6
+ 34 0.8 1.625
+ 34 0.8 1.65
+ 34 0.8 1.675
+ 34 0.8 1.7
+ 34 0.8 1.725
+ 34 0.8 1.75
+ 34 0.8 1.775
+ 34 0.8 1.8
+ 34 0.8 1.825
+ 34 0.8 1.85
+ 34 0.8 1.875
+ 34 0.8 1.9
+ 34 0.8 1.925
+ 34 0.8 1.95
+ 34 0.8 1.975
+ 34 0.8 2.0
+ 34 0.8 2.025
+ 34 0.8 2.05
+ 34 0.8 2.075
+ 34 0.8 2.1
+ 34 0.8 2.125
+ 34 0.8 2.15
+ 34 0.8 2.175
+ 34 0.8 2.2
+ 34 0.8 2.225
+ 34 0.8 2.25
+ 34 0.8 2.275
+ 34 0.8 2.3
+ 34 0.8 2.325
+ 34 0.8 2.35
+ 34 0.8 2.375
+ 34 0.8 2.4
+ 34 0.8 2.425
+ 34 0.8 2.45
+ 34 0.8 2.475
+ 34 0.8 2.5
+ 36 0.8 1.25
+ 36 0.8 1.275
+ 36 0.8 1.3
+ 36 0.8 1.325
+ 36 0.8 1.35
+ 36 0.8 1.375
+ 36 0.8 1.4
+ 36 0.8 1.425
+ 36 0.8 1.45
+ 36 0.8 1.475
+ 36 0.8 1.5
+ 36 0.8 1.525
+ 36 0.8 1.55
+ 36 0.8 1.575
+ 36 0.8 1.6
+ 36 0.8 1.625
+ 36 0.8 1.65
+ 36 0.8 1.675
+ 36 0.8 1.7
+ 36 0.8 1.725
+ 36 0.8 1.75
+ 36 0.8 1.775
+ 36 0.8 1.8
+ 36 0.8 1.825
+ 36 0.8 1.85
+ 36 0.8 1.875
+ 36 0.8 1.9
+ 36 0.8 1.925
+ 36 0.8 1.95
+ 36 0.8 1.975
+ 36 0.8 2.0
+ 36 0.8 2.025
+ 36 0.8 2.05
+ 36 0.8 2.075
+ 36 0.8 2.1
+ 36 0.8 2.125
+ 36 0.8 2.15
+ 36 0.8 2.175
+ 36 0.8 2.2
+ 36 0.8 2.225
+ 36 0.8 2.25
+ 36 0.8 2.275
+ 36 0.8 2.3
+ 36 0.8 2.325
+ 36 0.8 2.35
+ 36 0.8 2.375
+ 36 0.8 2.4
+ 36 0.8 2.425
+ 36 0.8 2.45
+ 36 0.8 2.475
+ 36 0.8 2.5
+ 38 0.8 1.25
+ 38 0.8 1.275
+ 38 0.8 1.3
+ 38 0.8 1.325
+ 38 0.8 1.35
+ 38 0.8 1.375
+ 38 0.8 1.4
+ 38 0.8 1.425
+ 38 0.8 1.45
+ 38 0.8 1.475
+ 38 0.8 1.5
+ 38 0.8 1.525
+ 38 0.8 1.55
+ 38 0.8 1.575
+ 38 0.8 1.6
+ 38 0.8 1.625
+ 38 0.8 1.65
+ 38 0.8 1.675
+ 38 0.8 1.7
+ 38 0.8 1.725
+ 38 0.8 1.75
+ 38 0.8 1.775
+ 38 0.8 1.8
+ 38 0.8 1.825
+ 38 0.8 1.85
+ 38 0.8 1.875
+ 38 0.8 1.9
+ 38 0.8 1.925
+ 38 0.8 1.95
+ 38 0.8 1.975
+ 38 0.8 2.0
+ 38 0.8 2.025
+ 38 0.8 2.05
+ 38 0.8 2.075
+ 38 0.8 2.1
+ 38 0.8 2.125
+ 38 0.8 2.15
+ 38 0.8 2.175
+ 38 0.8 2.2
+ 38 0.8 2.225
+ 38 0.8 2.25
+ 38 0.8 2.275
+ 38 0.8 2.3
+ 38 0.8 2.325
+ 38 0.8 2.35
+ 38 0.8 2.375
+ 38 0.8 2.4
+ 38 0.8 2.425
+ 38 0.8 2.45
+ 38 0.8 2.475
+ 38 0.8 2.5
+ 40 0.8 1.25
+ 40 0.8 1.275
+ 40 0.8 1.3
+ 40 0.8 1.325
+ 40 0.8 1.35
+ 40 0.8 1.375
+ 40 0.8 1.4
+ 40 0.8 1.425
+ 40 0.8 1.45
+ 40 0.8 1.475
+ 40 0.8 1.5
+ 40 0.8 1.525
+ 40 0.8 1.55
+ 40 0.8 1.575
+ 40 0.8 1.6
+ 40 0.8 1.625
+ 40 0.8 1.65
+ 40 0.8 1.675
+ 40 0.8 1.7
+ 40 0.8 1.725
+ 40 0.8 1.75
+ 40 0.8 1.775
+ 40 0.8 1.8
+ 40 0.8 1.825
+ 40 0.8 1.85
+ 40 0.8 1.875
+ 40 0.8 1.9
+ 40 0.8 1.925
+ 40 0.8 1.95
+ 40 0.8 1.975
+ 40 0.8 2.0
+ 40 0.8 2.025
+ 40 0.8 2.05
+ 40 0.8 2.075
+ 40 0.8 2.1
+ 40 0.8 2.125
+ 40 0.8 2.15
+ 40 0.8 2.175
+ 40 0.8 2.2
+ 40 0.8 2.225
+ 40 0.8 2.25
+ 40 0.8 2.275
+ 40 0.8 2.3
+ 40 0.8 2.325
+ 40 0.8 2.35
+ 40 0.8 2.375
+ 40 0.8 2.4
+ 40 0.8 2.425
+ 40 0.8 2.45
+ 40 0.8 2.475
+ 40 0.8 2.5
+ 42 0.8 1.25
+ 42 0.8 1.275
+ 42 0.8 1.3
+ 42 0.8 1.325
+ 42 0.8 1.35
+ 42 0.8 1.375
+ 42 0.8 1.4
+ 42 0.8 1.425
+ 42 0.8 1.45
+ 42 0.8 1.475
+ 42 0.8 1.5
+ 42 0.8 1.525
+ 42 0.8 1.55
+ 42 0.8 1.575
+ 42 0.8 1.6
+ 42 0.8 1.625
+ 42 0.8 1.65
+ 42 0.8 1.675
+ 42 0.8 1.7
+ 42 0.8 1.725
+ 42 0.8 1.75
+ 42 0.8 1.775
+ 42 0.8 1.8
+ 42 0.8 1.825
+ 42 0.8 1.85
+ 42 0.8 1.875
+ 42 0.8 1.9
+ 42 0.8 1.925
+ 42 0.8 1.95
+ 42 0.8 1.975
+ 42 0.8 2.0
+ 42 0.8 2.025
+ 42 0.8 2.05
+ 42 0.8 2.075
+ 42 0.8 2.1
+ 42 0.8 2.125
+ 42 0.8 2.15
+ 42 0.8 2.175
+ 42 0.8 2.2
+ 42 0.8 2.225
+ 42 0.8 2.25
+ 42 0.8 2.275
+ 42 0.8 2.3
+ 42 0.8 2.325
+ 42 0.8 2.35
+ 42 0.8 2.375
+ 42 0.8 2.4
+ 42 0.8 2.425
+ 42 0.8 2.45
+ 42 0.8 2.475
+ 42 0.8 2.5
+ 44 0.8 1.25
+ 44 0.8 1.275
+ 44 0.8 1.3
+ 44 0.8 1.325
+ 44 0.8 1.35
+ 44 0.8 1.375
+ 44 0.8 1.4
+ 44 0.8 1.425
+ 44 0.8 1.45
+ 44 0.8 1.475
+ 44 0.8 1.5
+ 44 0.8 1.525
+ 44 0.8 1.55
+ 44 0.8 1.575
+ 44 0.8 1.6
+ 44 0.8 1.625
+ 44 0.8 1.65
+ 44 0.8 1.675
+ 44 0.8 1.7
+ 44 0.8 1.725
+ 44 0.8 1.75
+ 44 0.8 1.775
+ 44 0.8 1.8
+ 44 0.8 1.825
+ 44 0.8 1.85
+ 44 0.8 1.875
+ 44 0.8 1.9
+ 44 0.8 1.925
+ 44 0.8 1.95
+ 44 0.8 1.975
+ 44 0.8 2.0
+ 44 0.8 2.025
+ 44 0.8 2.05
+ 44 0.8 2.075
+ 44 0.8 2.1
+ 44 0.8 2.125
+ 44 0.8 2.15
+ 44 0.8 2.175
+ 44 0.8 2.2
+ 44 0.8 2.225
+ 44 0.8 2.25
+ 44 0.8 2.275
+ 44 0.8 2.3
+ 44 0.8 2.325
+ 44 0.8 2.35
+ 44 0.8 2.375
+ 44 0.8 2.4
+ 44 0.8 2.425
+ 44 0.8 2.45
+ 44 0.8 2.475
+ 44 0.8 2.5
+ 46 0.8 1.25
+ 46 0.8 1.275
+ 46 0.8 1.3
+ 46 0.8 1.325
+ 46 0.8 1.35
+ 46 0.8 1.375
+ 46 0.8 1.4
+ 46 0.8 1.425
+ 46 0.8 1.45
+ 46 0.8 1.475
+ 46 0.8 1.5
+ 46 0.8 1.525
+ 46 0.8 1.55
+ 46 0.8 1.575
+ 46 0.8 1.6
+ 46 0.8 1.625
+ 46 0.8 1.65
+ 46 0.8 1.675
+ 46 0.8 1.7
+ 46 0.8 1.725
+ 46 0.8 1.75
+ 46 0.8 1.775
+ 46 0.8 1.8
+ 46 0.8 1.825
+ 46 0.8 1.85
+ 46 0.8 1.875
+ 46 0.8 1.9
+ 46 0.8 1.925
+ 46 0.8 1.95
+ 46 0.8 1.975
+ 46 0.8 2.0
+ 46 0.8 2.025
+ 46 0.8 2.05
+ 46 0.8 2.075
+ 46 0.8 2.1
+ 46 0.8 2.125
+ 46 0.8 2.15
+ 46 0.8 2.175
+ 46 0.8 2.2
+ 46 0.8 2.225
+ 46 0.8 2.25
+ 46 0.8 2.275
+ 46 0.8 2.3
+ 46 0.8 2.325
+ 46 0.8 2.35
+ 46 0.8 2.375
+ 46 0.8 2.4
+ 46 0.8 2.425
+ 46 0.8 2.45
+ 46 0.8 2.475
+ 46 0.8 2.5
+ 48 0.8 1.25
+ 48 0.8 1.275
+ 48 0.8 1.3
+ 48 0.8 1.325
+ 48 0.8 1.35
+ 48 0.8 1.375
+ 48 0.8 1.4
+ 48 0.8 1.425
+ 48 0.8 1.45
+ 48 0.8 1.475
+ 48 0.8 1.5
+ 48 0.8 1.525
+ 48 0.8 1.55
+ 48 0.8 1.575
+ 48 0.8 1.6
+ 48 0.8 1.625
+ 48 0.8 1.65
+ 48 0.8 1.675
+ 48 0.8 1.7
+ 48 0.8 1.725
+ 48 0.8 1.75
+ 48 0.8 1.775
+ 48 0.8 1.8
+ 48 0.8 1.825
+ 48 0.8 1.85
+ 48 0.8 1.875
+ 48 0.8 1.9
+ 48 0.8 1.925
+ 48 0.8 1.95
+ 48 0.8 1.975
+ 48 0.8 2.0
+ 48 0.8 2.025
+ 48 0.8 2.05
+ 48 0.8 2.075
+ 48 0.8 2.1
+ 48 0.8 2.125
+ 48 0.8 2.15
+ 48 0.8 2.175
+ 48 0.8 2.2
+ 48 0.8 2.225
+ 48 0.8 2.25
+ 48 0.8 2.275
+ 48 0.8 2.3
+ 48 0.8 2.325
+ 48 0.8 2.35
+ 48 0.8 2.375
+ 48 0.8 2.4
+ 48 0.8 2.425
+ 48 0.8 2.45
+ 48 0.8 2.475
+ 48 0.8 2.5
+ 50 0.8 1.25
+ 50 0.8 1.275
+ 50 0.8 1.3
+ 50 0.8 1.325
+ 50 0.8 1.35
+ 50 0.8 1.375
+ 50 0.8 1.4
+ 50 0.8 1.425
+ 50 0.8 1.45
+ 50 0.8 1.475
+ 50 0.8 1.5
+ 50 0.8 1.525
+ 50 0.8 1.55
+ 50 0.8 1.575
+ 50 0.8 1.6
+ 50 0.8 1.625
+ 50 0.8 1.65
+ 50 0.8 1.675
+ 50 0.8 1.7
+ 50 0.8 1.725
+ 50 0.8 1.75
+ 50 0.8 1.775
+ 50 0.8 1.8
+ 50 0.8 1.825
+ 50 0.8 1.85
+ 50 0.8 1.875
+ 50 0.8 1.9
+ 50 0.8 1.925
+ 50 0.8 1.95
+ 50 0.8 1.975
+ 50 0.8 2.0
+ 50 0.8 2.025
+ 50 0.8 2.05
+ 50 0.8 2.075
+ 50 0.8 2.1
+ 50 0.8 2.125
+ 50 0.8 2.15
+ 50 0.8 2.175
+ 50 0.8 2.2
+ 50 0.8 2.225
+ 50 0.8 2.25
+ 50 0.8 2.275
+ 50 0.8 2.3
+ 50 0.8 2.325
+ 50 0.8 2.35
+ 50 0.8 2.375
+ 50 0.8 2.4
+ 50 0.8 2.425
+ 50 0.8 2.45
+ 50 0.8 2.475
+ 50 0.8 2.5
+ 52 0.8 1.25
+ 52 0.8 1.275
+ 52 0.8 1.3
+ 52 0.8 1.325
+ 52 0.8 1.35
+ 52 0.8 1.375
+ 52 0.8 1.4
+ 52 0.8 1.425
+ 52 0.8 1.45
+ 52 0.8 1.475
+ 52 0.8 1.5
+ 52 0.8 1.525
+ 52 0.8 1.55
+ 52 0.8 1.575
+ 52 0.8 1.6
+ 52 0.8 1.625
+ 52 0.8 1.65
+ 52 0.8 1.675
+ 52 0.8 1.7
+ 52 0.8 1.725
+ 52 0.8 1.75
+ 52 0.8 1.775
+ 52 0.8 1.8
+ 52 0.8 1.825
+ 52 0.8 1.85
+ 52 0.8 1.875
+ 52 0.8 1.9
+ 52 0.8 1.925
+ 52 0.8 1.95
+ 52 0.8 1.975
+ 52 0.8 2.0
+ 52 0.8 2.025
+ 52 0.8 2.05
+ 52 0.8 2.075
+ 52 0.8 2.1
+ 52 0.8 2.125
+ 52 0.8 2.15
+ 52 0.8 2.175
+ 52 0.8 2.2
+ 52 0.8 2.225
+ 52 0.8 2.25
+ 52 0.8 2.275
+ 52 0.8 2.3
+ 52 0.8 2.325
+ 52 0.8 2.35
+ 52 0.8 2.375
+ 52 0.8 2.4
+ 52 0.8 2.425
+ 52 0.8 2.45
+ 52 0.8 2.475
+ 52 0.8 2.5
+ 54 0.8 1.25
+ 54 0.8 1.275
+ 54 0.8 1.3
+ 54 0.8 1.325
+ 54 0.8 1.35
+ 54 0.8 1.375
+ 54 0.8 1.4
+ 54 0.8 1.425
+ 54 0.8 1.45
+ 54 0.8 1.475
+ 54 0.8 1.5
+ 54 0.8 1.525
+ 54 0.8 1.55
+ 54 0.8 1.575
+ 54 0.8 1.6
+ 54 0.8 1.625
+ 54 0.8 1.65
+ 54 0.8 1.675
+ 54 0.8 1.7
+ 54 0.8 1.725
+ 54 0.8 1.75
+ 54 0.8 1.775
+ 54 0.8 1.8
+ 54 0.8 1.825
+ 54 0.8 1.85
+ 54 0.8 1.875
+ 54 0.8 1.9
+ 54 0.8 1.925
+ 54 0.8 1.95
+ 54 0.8 1.975
+ 54 0.8 2.0
+ 54 0.8 2.025
+ 54 0.8 2.05
+ 54 0.8 2.075
+ 54 0.8 2.1
+ 54 0.8 2.125
+ 54 0.8 2.15
+ 54 0.8 2.175
+ 54 0.8 2.2
+ 54 0.8 2.225
+ 54 0.8 2.25
+ 54 0.8 2.275
+ 54 0.8 2.3
+ 54 0.8 2.325
+ 54 0.8 2.35
+ 54 0.8 2.375
+ 54 0.8 2.4
+ 54 0.8 2.425
+ 54 0.8 2.45
+ 54 0.8 2.475
+ 54 0.8 2.5
+ 56 0.8 1.25
+ 56 0.8 1.275
+ 56 0.8 1.3
+ 56 0.8 1.325
+ 56 0.8 1.35
+ 56 0.8 1.375
+ 56 0.8 1.4
+ 56 0.8 1.425
+ 56 0.8 1.45
+ 56 0.8 1.475
+ 56 0.8 1.5
+ 56 0.8 1.525
+ 56 0.8 1.55
+ 56 0.8 1.575
+ 56 0.8 1.6
+ 56 0.8 1.625
+ 56 0.8 1.65
+ 56 0.8 1.675
+ 56 0.8 1.7
+ 56 0.8 1.725
+ 56 0.8 1.75
+ 56 0.8 1.775
+ 56 0.8 1.8
+ 56 0.8 1.825
+ 56 0.8 1.85
+ 56 0.8 1.875
+ 56 0.8 1.9
+ 56 0.8 1.925
+ 56 0.8 1.95
+ 56 0.8 1.975
+ 56 0.8 2.0
+ 56 0.8 2.025
+ 56 0.8 2.05
+ 56 0.8 2.075
+ 56 0.8 2.1
+ 56 0.8 2.125
+ 56 0.8 2.15
+ 56 0.8 2.175
+ 56 0.8 2.2
+ 56 0.8 2.225
+ 56 0.8 2.25
+ 56 0.8 2.275
+ 56 0.8 2.3
+ 56 0.8 2.325
+ 56 0.8 2.35
+ 56 0.8 2.375
+ 56 0.8 2.4
+ 56 0.8 2.425
+ 56 0.8 2.45
+ 56 0.8 2.475
+ 56 0.8 2.5
+ 58 0.8 1.25
+ 58 0.8 1.275
+ 58 0.8 1.3
+ 58 0.8 1.325
+ 58 0.8 1.35
+ 58 0.8 1.375
+ 58 0.8 1.4
+ 58 0.8 1.425
+ 58 0.8 1.45
+ 58 0.8 1.475
+ 58 0.8 1.5
+ 58 0.8 1.525
+ 58 0.8 1.55
+ 58 0.8 1.575
+ 58 0.8 1.6
+ 58 0.8 1.625
+ 58 0.8 1.65
+ 58 0.8 1.675
+ 58 0.8 1.7
+ 58 0.8 1.725
+ 58 0.8 1.75
+ 58 0.8 1.775
+ 58 0.8 1.8
+ 58 0.8 1.825
+ 58 0.8 1.85
+ 58 0.8 1.875
+ 58 0.8 1.9
+ 58 0.8 1.925
+ 58 0.8 1.95
+ 58 0.8 1.975
+ 58 0.8 2.0
+ 58 0.8 2.025
+ 58 0.8 2.05
+ 58 0.8 2.075
+ 58 0.8 2.1
+ 58 0.8 2.125
+ 58 0.8 2.15
+ 58 0.8 2.175
+ 58 0.8 2.2
+ 58 0.8 2.225
+ 58 0.8 2.25
+ 58 0.8 2.275
+ 58 0.8 2.3
+ 58 0.8 2.325
+ 58 0.8 2.35
+ 58 0.8 2.375
+ 58 0.8 2.4
+ 58 0.8 2.425
+ 58 0.8 2.45
+ 58 0.8 2.475
+ 58 0.8 2.5
+ 60 0.8 1.25
+ 60 0.8 1.275
+ 60 0.8 1.3
+ 60 0.8 1.325
+ 60 0.8 1.35
+ 60 0.8 1.375
+ 60 0.8 1.4
+ 60 0.8 1.425
+ 60 0.8 1.45
+ 60 0.8 1.475
+ 60 0.8 1.5
+ 60 0.8 1.525
+ 60 0.8 1.55
+ 60 0.8 1.575
+ 60 0.8 1.6
+ 60 0.8 1.625
+ 60 0.8 1.65
+ 60 0.8 1.675
+ 60 0.8 1.7
+ 60 0.8 1.725
+ 60 0.8 1.75
+ 60 0.8 1.775
+ 60 0.8 1.8
+ 60 0.8 1.825
+ 60 0.8 1.85
+ 60 0.8 1.875
+ 60 0.8 1.9
+ 60 0.8 1.925
+ 60 0.8 1.95
+ 60 0.8 1.975
+ 60 0.8 2.0
+ 60 0.8 2.025
+ 60 0.8 2.05
+ 60 0.8 2.075
+ 60 0.8 2.1
+ 60 0.8 2.125
+ 60 0.8 2.15
+ 60 0.8 2.175
+ 60 0.8 2.2
+ 60 0.8 2.225
+ 60 0.8 2.25
+ 60 0.8 2.275
+ 60 0.8 2.3
+ 60 0.8 2.325
+ 60 0.8 2.35
+ 60 0.8 2.375
+ 60 0.8 2.4
+ 60 0.8 2.425
+ 60 0.8 2.45
+ 60 0.8 2.475
+ 60 0.8 2.5
+ 62 0.8 1.25
+ 62 0.8 1.275
+ 62 0.8 1.3
+ 62 0.8 1.325
+ 62 0.8 1.35
+ 62 0.8 1.375
+ 62 0.8 1.4
+ 62 0.8 1.425
+ 62 0.8 1.45
+ 62 0.8 1.475
+ 62 0.8 1.5
+ 62 0.8 1.525
+ 62 0.8 1.55
+ 62 0.8 1.575
+ 62 0.8 1.6
+ 62 0.8 1.625
+ 62 0.8 1.65
+ 62 0.8 1.675
+ 62 0.8 1.7
+ 62 0.8 1.725
+ 62 0.8 1.75
+ 62 0.8 1.775
+ 62 0.8 1.8
+ 62 0.8 1.825
+ 62 0.8 1.85
+ 62 0.8 1.875
+ 62 0.8 1.9
+ 62 0.8 1.925
+ 62 0.8 1.95
+ 62 0.8 1.975
+ 62 0.8 2.0
+ 62 0.8 2.025
+ 62 0.8 2.05
+ 62 0.8 2.075
+ 62 0.8 2.1
+ 62 0.8 2.125
+ 62 0.8 2.15
+ 62 0.8 2.175
+ 62 0.8 2.2
+ 62 0.8 2.225
+ 62 0.8 2.25
+ 62 0.8 2.275
+ 62 0.8 2.3
+ 62 0.8 2.325
+ 62 0.8 2.35
+ 62 0.8 2.375
+ 62 0.8 2.4
+ 62 0.8 2.425
+ 62 0.8 2.45
+ 62 0.8 2.475
+ 62 0.8 2.5
+ 64 0.8 1.25
+ 64 0.8 1.275
+ 64 0.8 1.3
+ 64 0.8 1.325
+ 64 0.8 1.35
+ 64 0.8 1.375
+ 64 0.8 1.4
+ 64 0.8 1.425
+ 64 0.8 1.45
+ 64 0.8 1.475
+ 64 0.8 1.5
+ 64 0.8 1.525
+ 64 0.8 1.55
+ 64 0.8 1.575
+ 64 0.8 1.6
+ 64 0.8 1.625
+ 64 0.8 1.65
+ 64 0.8 1.675
+ 64 0.8 1.7
+ 64 0.8 1.725
+ 64 0.8 1.75
+ 64 0.8 1.775
+ 64 0.8 1.8
+ 64 0.8 1.825
+ 64 0.8 1.85
+ 64 0.8 1.875
+ 64 0.8 1.9
+ 64 0.8 1.925
+ 64 0.8 1.95
+ 64 0.8 1.975
+ 64 0.8 2.0
+ 64 0.8 2.025
+ 64 0.8 2.05
+ 64 0.8 2.075
+ 64 0.8 2.1
+ 64 0.8 2.125
+ 64 0.8 2.15
+ 64 0.8 2.175
+ 64 0.8 2.2
+ 64 0.8 2.225
+ 64 0.8 2.25
+ 64 0.8 2.275
+ 64 0.8 2.3
+ 64 0.8 2.325
+ 64 0.8 2.35
+ 64 0.8 2.375
+ 64 0.8 2.4
+ 64 0.8 2.425
+ 64 0.8 2.45
+ 64 0.8 2.475
+ 64 0.8 2.5
+ 66 0.8 1.25
+ 66 0.8 1.275
+ 66 0.8 1.3
+ 66 0.8 1.325
+ 66 0.8 1.35
+ 66 0.8 1.375
+ 66 0.8 1.4
+ 66 0.8 1.425
+ 66 0.8 1.45
+ 66 0.8 1.475
+ 66 0.8 1.5
+ 66 0.8 1.525
+ 66 0.8 1.55
+ 66 0.8 1.575
+ 66 0.8 1.6
+ 66 0.8 1.625
+ 66 0.8 1.65
+ 66 0.8 1.675
+ 66 0.8 1.7
+ 66 0.8 1.725
+ 66 0.8 1.75
+ 66 0.8 1.775
+ 66 0.8 1.8
+ 66 0.8 1.825
+ 66 0.8 1.85
+ 66 0.8 1.875
+ 66 0.8 1.9
+ 66 0.8 1.925
+ 66 0.8 1.95
+ 66 0.8 1.975
+ 66 0.8 2.0
+ 66 0.8 2.025
+ 66 0.8 2.05
+ 66 0.8 2.075
+ 66 0.8 2.1
+ 66 0.8 2.125
+ 66 0.8 2.15
+ 66 0.8 2.175
+ 66 0.8 2.2
+ 66 0.8 2.225
+ 66 0.8 2.25
+ 66 0.8 2.275
+ 66 0.8 2.3
+ 66 0.8 2.325
+ 66 0.8 2.35
+ 66 0.8 2.375
+ 66 0.8 2.4
+ 66 0.8 2.425
+ 66 0.8 2.45
+ 66 0.8 2.475
+ 66 0.8 2.5
+ 68 0.8 1.25
+ 68 0.8 1.275
+ 68 0.8 1.3
+ 68 0.8 1.325
+ 68 0.8 1.35
+ 68 0.8 1.375
+ 68 0.8 1.4
+ 68 0.8 1.425
+ 68 0.8 1.45
+ 68 0.8 1.475
+ 68 0.8 1.5
+ 68 0.8 1.525
+ 68 0.8 1.55
+ 68 0.8 1.575
+ 68 0.8 1.6
+ 68 0.8 1.625
+ 68 0.8 1.65
+ 68 0.8 1.675
+ 68 0.8 1.7
+ 68 0.8 1.725
+ 68 0.8 1.75
+ 68 0.8 1.775
+ 68 0.8 1.8
+ 68 0.8 1.825
+ 68 0.8 1.85
+ 68 0.8 1.875
+ 68 0.8 1.9
+ 68 0.8 1.925
+ 68 0.8 1.95
+ 68 0.8 1.975
+ 68 0.8 2.0
+ 68 0.8 2.025
+ 68 0.8 2.05
+ 68 0.8 2.075
+ 68 0.8 2.1
+ 68 0.8 2.125
+ 68 0.8 2.15
+ 68 0.8 2.175
+ 68 0.8 2.2
+ 68 0.8 2.225
+ 68 0.8 2.25
+ 68 0.8 2.275
+ 68 0.8 2.3
+ 68 0.8 2.325
+ 68 0.8 2.35
+ 68 0.8 2.375
+ 68 0.8 2.4
+ 68 0.8 2.425
+ 68 0.8 2.45
+ 68 0.8 2.475
+ 68 0.8 2.5
+ 70 0.8 1.25
+ 70 0.8 1.275
+ 70 0.8 1.3
+ 70 0.8 1.325
+ 70 0.8 1.35
+ 70 0.8 1.375
+ 70 0.8 1.4
+ 70 0.8 1.425
+ 70 0.8 1.45
+ 70 0.8 1.475
+ 70 0.8 1.5
+ 70 0.8 1.525
+ 70 0.8 1.55
+ 70 0.8 1.575
+ 70 0.8 1.6
+ 70 0.8 1.625
+ 70 0.8 1.65
+ 70 0.8 1.675
+ 70 0.8 1.7
+ 70 0.8 1.725
+ 70 0.8 1.75
+ 70 0.8 1.775
+ 70 0.8 1.8
+ 70 0.8 1.825
+ 70 0.8 1.85
+ 70 0.8 1.875
+ 70 0.8 1.9
+ 70 0.8 1.925
+ 70 0.8 1.95
+ 70 0.8 1.975
+ 70 0.8 2.0
+ 70 0.8 2.025
+ 70 0.8 2.05
+ 70 0.8 2.075
+ 70 0.8 2.1
+ 70 0.8 2.125
+ 70 0.8 2.15
+ 70 0.8 2.175
+ 70 0.8 2.2
+ 70 0.8 2.225
+ 70 0.8 2.25
+ 70 0.8 2.275
+ 70 0.8 2.3
+ 70 0.8 2.325
+ 70 0.8 2.35
+ 70 0.8 2.375
+ 70 0.8 2.4
+ 70 0.8 2.425
+ 70 0.8 2.45
+ 70 0.8 2.475
+ 70 0.8 2.5
+ 72 0.8 1.25
+ 72 0.8 1.275
+ 72 0.8 1.3
+ 72 0.8 1.325
+ 72 0.8 1.35
+ 72 0.8 1.375
+ 72 0.8 1.4
+ 72 0.8 1.425
+ 72 0.8 1.45
+ 72 0.8 1.475
+ 72 0.8 1.5
+ 72 0.8 1.525
+ 72 0.8 1.55
+ 72 0.8 1.575
+ 72 0.8 1.6
+ 72 0.8 1.625
+ 72 0.8 1.65
+ 72 0.8 1.675
+ 72 0.8 1.7
+ 72 0.8 1.725
+ 72 0.8 1.75
+ 72 0.8 1.775
+ 72 0.8 1.8
+ 72 0.8 1.825
+ 72 0.8 1.85
+ 72 0.8 1.875
+ 72 0.8 1.9
+ 72 0.8 1.925
+ 72 0.8 1.95
+ 72 0.8 1.975
+ 72 0.8 2.0
+ 72 0.8 2.025
+ 72 0.8 2.05
+ 72 0.8 2.075
+ 72 0.8 2.1
+ 72 0.8 2.125
+ 72 0.8 2.15
+ 72 0.8 2.175
+ 72 0.8 2.2
+ 72 0.8 2.225
+ 72 0.8 2.25
+ 72 0.8 2.275
+ 72 0.8 2.3
+ 72 0.8 2.325
+ 72 0.8 2.35
+ 72 0.8 2.375
+ 72 0.8 2.4
+ 72 0.8 2.425
+ 72 0.8 2.45
+ 72 0.8 2.475
+ 72 0.8 2.5
+ 74 0.8 1.25
+ 74 0.8 1.275
+ 74 0.8 1.3
+ 74 0.8 1.325
+ 74 0.8 1.35
+ 74 0.8 1.375
+ 74 0.8 1.4
+ 74 0.8 1.425
+ 74 0.8 1.45
+ 74 0.8 1.475
+ 74 0.8 1.5
+ 74 0.8 1.525
+ 74 0.8 1.55
+ 74 0.8 1.575
+ 74 0.8 1.6
+ 74 0.8 1.625
+ 74 0.8 1.65
+ 74 0.8 1.675
+ 74 0.8 1.7
+ 74 0.8 1.725
+ 74 0.8 1.75
+ 74 0.8 1.775
+ 74 0.8 1.8
+ 74 0.8 1.825
+ 74 0.8 1.85
+ 74 0.8 1.875
+ 74 0.8 1.9
+ 74 0.8 1.925
+ 74 0.8 1.95
+ 74 0.8 1.975
+ 74 0.8 2.0
+ 74 0.8 2.025
+ 74 0.8 2.05
+ 74 0.8 2.075
+ 74 0.8 2.1
+ 74 0.8 2.125
+ 74 0.8 2.15
+ 74 0.8 2.175
+ 74 0.8 2.2
+ 74 0.8 2.225
+ 74 0.8 2.25
+ 74 0.8 2.275
+ 74 0.8 2.3
+ 74 0.8 2.325
+ 74 0.8 2.35
+ 74 0.8 2.375
+ 74 0.8 2.4
+ 74 0.8 2.425
+ 74 0.8 2.45
+ 74 0.8 2.475
+ 74 0.8 2.5
+ 76 0.8 1.25
+ 76 0.8 1.275
+ 76 0.8 1.3
+ 76 0.8 1.325
+ 76 0.8 1.35
+ 76 0.8 1.375
+ 76 0.8 1.4
+ 76 0.8 1.425
+ 76 0.8 1.45
+ 76 0.8 1.475
+ 76 0.8 1.5
+ 76 0.8 1.525
+ 76 0.8 1.55
+ 76 0.8 1.575
+ 76 0.8 1.6
+ 76 0.8 1.625
+ 76 0.8 1.65
+ 76 0.8 1.675
+ 76 0.8 1.7
+ 76 0.8 1.725
+ 76 0.8 1.75
+ 76 0.8 1.775
+ 76 0.8 1.8
+ 76 0.8 1.825
+ 76 0.8 1.85
+ 76 0.8 1.875
+ 76 0.8 1.9
+ 76 0.8 1.925
+ 76 0.8 1.95
+ 76 0.8 1.975
+ 76 0.8 2.0
+ 76 0.8 2.025
+ 76 0.8 2.05
+ 76 0.8 2.075
+ 76 0.8 2.1
+ 76 0.8 2.125
+ 76 0.8 2.15
+ 76 0.8 2.175
+ 76 0.8 2.2
+ 76 0.8 2.225
+ 76 0.8 2.25
+ 76 0.8 2.275
+ 76 0.8 2.3
+ 76 0.8 2.325
+ 76 0.8 2.35
+ 76 0.8 2.375
+ 76 0.8 2.4
+ 76 0.8 2.425
+ 76 0.8 2.45
+ 76 0.8 2.475
+ 76 0.8 2.5
+ 78 0.8 1.25
+ 78 0.8 1.275
+ 78 0.8 1.3
+ 78 0.8 1.325
+ 78 0.8 1.35
+ 78 0.8 1.375
+ 78 0.8 1.4
+ 78 0.8 1.425
+ 78 0.8 1.45
+ 78 0.8 1.475
+ 78 0.8 1.5
+ 78 0.8 1.525
+ 78 0.8 1.55
+ 78 0.8 1.575
+ 78 0.8 1.6
+ 78 0.8 1.625
+ 78 0.8 1.65
+ 78 0.8 1.675
+ 78 0.8 1.7
+ 78 0.8 1.725
+ 78 0.8 1.75
+ 78 0.8 1.775
+ 78 0.8 1.8
+ 78 0.8 1.825
+ 78 0.8 1.85
+ 78 0.8 1.875
+ 78 0.8 1.9
+ 78 0.8 1.925
+ 78 0.8 1.95
+ 78 0.8 1.975
+ 78 0.8 2.0
+ 78 0.8 2.025
+ 78 0.8 2.05
+ 78 0.8 2.075
+ 78 0.8 2.1
+ 78 0.8 2.125
+ 78 0.8 2.15
+ 78 0.8 2.175
+ 78 0.8 2.2
+ 78 0.8 2.225
+ 78 0.8 2.25
+ 78 0.8 2.275
+ 78 0.8 2.3
+ 78 0.8 2.325
+ 78 0.8 2.35
+ 78 0.8 2.375
+ 78 0.8 2.4
+ 78 0.8 2.425
+ 78 0.8 2.45
+ 78 0.8 2.475
+ 78 0.8 2.5
+ 80 0.8 1.25
+ 80 0.8 1.275
+ 80 0.8 1.3
+ 80 0.8 1.325
+ 80 0.8 1.35
+ 80 0.8 1.375
+ 80 0.8 1.4
+ 80 0.8 1.425
+ 80 0.8 1.45
+ 80 0.8 1.475
+ 80 0.8 1.5
+ 80 0.8 1.525
+ 80 0.8 1.55
+ 80 0.8 1.575
+ 80 0.8 1.6
+ 80 0.8 1.625
+ 80 0.8 1.65
+ 80 0.8 1.675
+ 80 0.8 1.7
+ 80 0.8 1.725
+ 80 0.8 1.75
+ 80 0.8 1.775
+ 80 0.8 1.8
+ 80 0.8 1.825
+ 80 0.8 1.85
+ 80 0.8 1.875
+ 80 0.8 1.9
+ 80 0.8 1.925
+ 80 0.8 1.95
+ 80 0.8 1.975
+ 80 0.8 2.0
+ 80 0.8 2.025
+ 80 0.8 2.05
+ 80 0.8 2.075
+ 80 0.8 2.1
+ 80 0.8 2.125
+ 80 0.8 2.15
+ 80 0.8 2.175
+ 80 0.8 2.2
+ 80 0.8 2.225
+ 80 0.8 2.25
+ 80 0.8 2.275
+ 80 0.8 2.3
+ 80 0.8 2.325
+ 80 0.8 2.35
+ 80 0.8 2.375
+ 80 0.8 2.4
+ 80 0.8 2.425
+ 80 0.8 2.45
+ 80 0.8 2.475
+ 80 0.8 2.5
+ 82 0.8 1.25
+ 82 0.8 1.275
+ 82 0.8 1.3
+ 82 0.8 1.325
+ 82 0.8 1.35
+ 82 0.8 1.375
+ 82 0.8 1.4
+ 82 0.8 1.425
+ 82 0.8 1.45
+ 82 0.8 1.475
+ 82 0.8 1.5
+ 82 0.8 1.525
+ 82 0.8 1.55
+ 82 0.8 1.575
+ 82 0.8 1.6
+ 82 0.8 1.625
+ 82 0.8 1.65
+ 82 0.8 1.675
+ 82 0.8 1.7
+ 82 0.8 1.725
+ 82 0.8 1.75
+ 82 0.8 1.775
+ 82 0.8 1.8
+ 82 0.8 1.825
+ 82 0.8 1.85
+ 82 0.8 1.875
+ 82 0.8 1.9
+ 82 0.8 1.925
+ 82 0.8 1.95
+ 82 0.8 1.975
+ 82 0.8 2.0
+ 82 0.8 2.025
+ 82 0.8 2.05
+ 82 0.8 2.075
+ 82 0.8 2.1
+ 82 0.8 2.125
+ 82 0.8 2.15
+ 82 0.8 2.175
+ 82 0.8 2.2
+ 82 0.8 2.225
+ 82 0.8 2.25
+ 82 0.8 2.275
+ 82 0.8 2.3
+ 82 0.8 2.325
+ 82 0.8 2.35
+ 82 0.8 2.375
+ 82 0.8 2.4
+ 82 0.8 2.425
+ 82 0.8 2.45
+ 82 0.8 2.475
+ 82 0.8 2.5
+ 84 0.8 1.25
+ 84 0.8 1.275
+ 84 0.8 1.3
+ 84 0.8 1.325
+ 84 0.8 1.35
+ 84 0.8 1.375
+ 84 0.8 1.4
+ 84 0.8 1.425
+ 84 0.8 1.45
+ 84 0.8 1.475
+ 84 0.8 1.5
+ 84 0.8 1.525
+ 84 0.8 1.55
+ 84 0.8 1.575
+ 84 0.8 1.6
+ 84 0.8 1.625
+ 84 0.8 1.65
+ 84 0.8 1.675
+ 84 0.8 1.7
+ 84 0.8 1.725
+ 84 0.8 1.75
+ 84 0.8 1.775
+ 84 0.8 1.8
+ 84 0.8 1.825
+ 84 0.8 1.85
+ 84 0.8 1.875
+ 84 0.8 1.9
+ 84 0.8 1.925
+ 84 0.8 1.95
+ 84 0.8 1.975
+ 84 0.8 2.0
+ 84 0.8 2.025
+ 84 0.8 2.05
+ 84 0.8 2.075
+ 84 0.8 2.1
+ 84 0.8 2.125
+ 84 0.8 2.15
+ 84 0.8 2.175
+ 84 0.8 2.2
+ 84 0.8 2.225
+ 84 0.8 2.25
+ 84 0.8 2.275
+ 84 0.8 2.3
+ 84 0.8 2.325
+ 84 0.8 2.35
+ 84 0.8 2.375
+ 84 0.8 2.4
+ 84 0.8 2.425
+ 84 0.8 2.45
+ 84 0.8 2.475
+ 84 0.8 2.5
+ 86 0.8 1.25
+ 86 0.8 1.275
+ 86 0.8 1.3
+ 86 0.8 1.325
+ 86 0.8 1.35
+ 86 0.8 1.375
+ 86 0.8 1.4
+ 86 0.8 1.425
+ 86 0.8 1.45
+ 86 0.8 1.475
+ 86 0.8 1.5
+ 86 0.8 1.525
+ 86 0.8 1.55
+ 86 0.8 1.575
+ 86 0.8 1.6
+ 86 0.8 1.625
+ 86 0.8 1.65
+ 86 0.8 1.675
+ 86 0.8 1.7
+ 86 0.8 1.725
+ 86 0.8 1.75
+ 86 0.8 1.775
+ 86 0.8 1.8
+ 86 0.8 1.825
+ 86 0.8 1.85
+ 86 0.8 1.875
+ 86 0.8 1.9
+ 86 0.8 1.925
+ 86 0.8 1.95
+ 86 0.8 1.975
+ 86 0.8 2.0
+ 86 0.8 2.025
+ 86 0.8 2.05
+ 86 0.8 2.075
+ 86 0.8 2.1
+ 86 0.8 2.125
+ 86 0.8 2.15
+ 86 0.8 2.175
+ 86 0.8 2.2
+ 86 0.8 2.225
+ 86 0.8 2.25
+ 86 0.8 2.275
+ 86 0.8 2.3
+ 86 0.8 2.325
+ 86 0.8 2.35
+ 86 0.8 2.375
+ 86 0.8 2.4
+ 86 0.8 2.425
+ 86 0.8 2.45
+ 86 0.8 2.475
+ 86 0.8 2.5
+ 88 0.8 1.25
+ 88 0.8 1.275
+ 88 0.8 1.3
+ 88 0.8 1.325
+ 88 0.8 1.35
+ 88 0.8 1.375
+ 88 0.8 1.4
+ 88 0.8 1.425
+ 88 0.8 1.45
+ 88 0.8 1.475
+ 88 0.8 1.5
+ 88 0.8 1.525
+ 88 0.8 1.55
+ 88 0.8 1.575
+ 88 0.8 1.6
+ 88 0.8 1.625
+ 88 0.8 1.65
+ 88 0.8 1.675
+ 88 0.8 1.7
+ 88 0.8 1.725
+ 88 0.8 1.75
+ 88 0.8 1.775
+ 88 0.8 1.8
+ 88 0.8 1.825
+ 88 0.8 1.85
+ 88 0.8 1.875
+ 88 0.8 1.9
+ 88 0.8 1.925
+ 88 0.8 1.95
+ 88 0.8 1.975
+ 88 0.8 2.0
+ 88 0.8 2.025
+ 88 0.8 2.05
+ 88 0.8 2.075
+ 88 0.8 2.1
+ 88 0.8 2.125
+ 88 0.8 2.15
+ 88 0.8 2.175
+ 88 0.8 2.2
+ 88 0.8 2.225
+ 88 0.8 2.25
+ 88 0.8 2.275
+ 88 0.8 2.3
+ 88 0.8 2.325
+ 88 0.8 2.35
+ 88 0.8 2.375
+ 88 0.8 2.4
+ 88 0.8 2.425
+ 88 0.8 2.45
+ 88 0.8 2.475
+ 88 0.8 2.5
+ 90 0.8 1.25
+ 90 0.8 1.275
+ 90 0.8 1.3
+ 90 0.8 1.325
+ 90 0.8 1.35
+ 90 0.8 1.375
+ 90 0.8 1.4
+ 90 0.8 1.425
+ 90 0.8 1.45
+ 90 0.8 1.475
+ 90 0.8 1.5
+ 90 0.8 1.525
+ 90 0.8 1.55
+ 90 0.8 1.575
+ 90 0.8 1.6
+ 90 0.8 1.625
+ 90 0.8 1.65
+ 90 0.8 1.675
+ 90 0.8 1.7
+ 90 0.8 1.725
+ 90 0.8 1.75
+ 90 0.8 1.775
+ 90 0.8 1.8
+ 90 0.8 1.825
+ 90 0.8 1.85
+ 90 0.8 1.875
+ 90 0.8 1.9
+ 90 0.8 1.925
+ 90 0.8 1.95
+ 90 0.8 1.975
+ 90 0.8 2.0
+ 90 0.8 2.025
+ 90 0.8 2.05
+ 90 0.8 2.075
+ 90 0.8 2.1
+ 90 0.8 2.125
+ 90 0.8 2.15
+ 90 0.8 2.175
+ 90 0.8 2.2
+ 90 0.8 2.225
+ 90 0.8 2.25
+ 90 0.8 2.275
+ 90 0.8 2.3
+ 90 0.8 2.325
+ 90 0.8 2.35
+ 90 0.8 2.375
+ 90 0.8 2.4
+ 90 0.8 2.425
+ 90 0.8 2.45
+ 90 0.8 2.475
+ 90 0.8 2.5
+ 92 0.8 1.25
+ 92 0.8 1.275
+ 92 0.8 1.3
+ 92 0.8 1.325
+ 92 0.8 1.35
+ 92 0.8 1.375
+ 92 0.8 1.4
+ 92 0.8 1.425
+ 92 0.8 1.45
+ 92 0.8 1.475
+ 92 0.8 1.5
+ 92 0.8 1.525
+ 92 0.8 1.55
+ 92 0.8 1.575
+ 92 0.8 1.6
+ 92 0.8 1.625
+ 92 0.8 1.65
+ 92 0.8 1.675
+ 92 0.8 1.7
+ 92 0.8 1.725
+ 92 0.8 1.75
+ 92 0.8 1.775
+ 92 0.8 1.8
+ 92 0.8 1.825
+ 92 0.8 1.85
+ 92 0.8 1.875
+ 92 0.8 1.9
+ 92 0.8 1.925
+ 92 0.8 1.95
+ 92 0.8 1.975
+ 92 0.8 2.0
+ 92 0.8 2.025
+ 92 0.8 2.05
+ 92 0.8 2.075
+ 92 0.8 2.1
+ 92 0.8 2.125
+ 92 0.8 2.15
+ 92 0.8 2.175
+ 92 0.8 2.2
+ 92 0.8 2.225
+ 92 0.8 2.25
+ 92 0.8 2.275
+ 92 0.8 2.3
+ 92 0.8 2.325
+ 92 0.8 2.35
+ 92 0.8 2.375
+ 92 0.8 2.4
+ 92 0.8 2.425
+ 92 0.8 2.45
+ 92 0.8 2.475
+ 92 0.8 2.5
+ 94 0.8 1.25
+ 94 0.8 1.275
+ 94 0.8 1.3
+ 94 0.8 1.325
+ 94 0.8 1.35
+ 94 0.8 1.375
+ 94 0.8 1.4
+ 94 0.8 1.425
+ 94 0.8 1.45
+ 94 0.8 1.475
+ 94 0.8 1.5
+ 94 0.8 1.525
+ 94 0.8 1.55
+ 94 0.8 1.575
+ 94 0.8 1.6
+ 94 0.8 1.625
+ 94 0.8 1.65
+ 94 0.8 1.675
+ 94 0.8 1.7
+ 94 0.8 1.725
+ 94 0.8 1.75
+ 94 0.8 1.775
+ 94 0.8 1.8
+ 94 0.8 1.825
+ 94 0.8 1.85
+ 94 0.8 1.875
+ 94 0.8 1.9
+ 94 0.8 1.925
+ 94 0.8 1.95
+ 94 0.8 1.975
+ 94 0.8 2.0
+ 94 0.8 2.025
+ 94 0.8 2.05
+ 94 0.8 2.075
+ 94 0.8 2.1
+ 94 0.8 2.125
+ 94 0.8 2.15
+ 94 0.8 2.175
+ 94 0.8 2.2
+ 94 0.8 2.225
+ 94 0.8 2.25
+ 94 0.8 2.275
+ 94 0.8 2.3
+ 94 0.8 2.325
+ 94 0.8 2.35
+ 94 0.8 2.375
+ 94 0.8 2.4
+ 94 0.8 2.425
+ 94 0.8 2.45
+ 94 0.8 2.475
+ 94 0.8 2.5
+ 96 0.8 1.25
+ 96 0.8 1.275
+ 96 0.8 1.3
+ 96 0.8 1.325
+ 96 0.8 1.35
+ 96 0.8 1.375
+ 96 0.8 1.4
+ 96 0.8 1.425
+ 96 0.8 1.45
+ 96 0.8 1.475
+ 96 0.8 1.5
+ 96 0.8 1.525
+ 96 0.8 1.55
+ 96 0.8 1.575
+ 96 0.8 1.6
+ 96 0.8 1.625
+ 96 0.8 1.65
+ 96 0.8 1.675
+ 96 0.8 1.7
+ 96 0.8 1.725
+ 96 0.8 1.75
+ 96 0.8 1.775
+ 96 0.8 1.8
+ 96 0.8 1.825
+ 96 0.8 1.85
+ 96 0.8 1.875
+ 96 0.8 1.9
+ 96 0.8 1.925
+ 96 0.8 1.95
+ 96 0.8 1.975
+ 96 0.8 2.0
+ 96 0.8 2.025
+ 96 0.8 2.05
+ 96 0.8 2.075
+ 96 0.8 2.1
+ 96 0.8 2.125
+ 96 0.8 2.15
+ 96 0.8 2.175
+ 96 0.8 2.2
+ 96 0.8 2.225
+ 96 0.8 2.25
+ 96 0.8 2.275
+ 96 0.8 2.3
+ 96 0.8 2.325
+ 96 0.8 2.35
+ 96 0.8 2.375
+ 96 0.8 2.4
+ 96 0.8 2.425
+ 96 0.8 2.45
+ 96 0.8 2.475
+ 96 0.8 2.5
+ 98 0.8 1.25
+ 98 0.8 1.275
+ 98 0.8 1.3
+ 98 0.8 1.325
+ 98 0.8 1.35
+ 98 0.8 1.375
+ 98 0.8 1.4
+ 98 0.8 1.425
+ 98 0.8 1.45
+ 98 0.8 1.475
+ 98 0.8 1.5
+ 98 0.8 1.525
+ 98 0.8 1.55
+ 98 0.8 1.575
+ 98 0.8 1.6
+ 98 0.8 1.625
+ 98 0.8 1.65
+ 98 0.8 1.675
+ 98 0.8 1.7
+ 98 0.8 1.725
+ 98 0.8 1.75
+ 98 0.8 1.775
+ 98 0.8 1.8
+ 98 0.8 1.825
+ 98 0.8 1.85
+ 98 0.8 1.875
+ 98 0.8 1.9
+ 98 0.8 1.925
+ 98 0.8 1.95
+ 98 0.8 1.975
+ 98 0.8 2.0
+ 98 0.8 2.025
+ 98 0.8 2.05
+ 98 0.8 2.075
+ 98 0.8 2.1
+ 98 0.8 2.125
+ 98 0.8 2.15
+ 98 0.8 2.175
+ 98 0.8 2.2
+ 98 0.8 2.225
+ 98 0.8 2.25
+ 98 0.8 2.275
+ 98 0.8 2.3
+ 98 0.8 2.325
+ 98 0.8 2.35
+ 98 0.8 2.375
+ 98 0.8 2.4
+ 98 0.8 2.425
+ 98 0.8 2.45
+ 98 0.8 2.475
+ 98 0.8 2.5
+ 100 0.8 1.25
+ 100 0.8 1.275
+ 100 0.8 1.3
+ 100 0.8 1.325
+ 100 0.8 1.35
+ 100 0.8 1.375
+ 100 0.8 1.4
+ 100 0.8 1.425
+ 100 0.8 1.45
+ 100 0.8 1.475
+ 100 0.8 1.5
+ 100 0.8 1.525
+ 100 0.8 1.55
+ 100 0.8 1.575
+ 100 0.8 1.6
+ 100 0.8 1.625
+ 100 0.8 1.65
+ 100 0.8 1.675
+ 100 0.8 1.7
+ 100 0.8 1.725
+ 100 0.8 1.75
+ 100 0.8 1.775
+ 100 0.8 1.8
+ 100 0.8 1.825
+ 100 0.8 1.85
+ 100 0.8 1.875
+ 100 0.8 1.9
+ 100 0.8 1.925
+ 100 0.8 1.95
+ 100 0.8 1.975
+ 100 0.8 2.0
+ 100 0.8 2.025
+ 100 0.8 2.05
+ 100 0.8 2.075
+ 100 0.8 2.1
+ 100 0.8 2.125
+ 100 0.8 2.15
+ 100 0.8 2.175
+ 100 0.8 2.2
+ 100 0.8 2.225
+ 100 0.8 2.25
+ 100 0.8 2.275
+ 100 0.8 2.3
+ 100 0.8 2.325
+ 100 0.8 2.35
+ 100 0.8 2.375
+ 100 0.8 2.4
+ 100 0.8 2.425
+ 100 0.8 2.45
+ 100 0.8 2.475
+ 100 0.8 2.5
.ENDDATA
