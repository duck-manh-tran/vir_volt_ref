
.option MEASFORM=3
.param vdd=0.8
.param vinit=0.4

.ic v(vp)='vinit+0.01'

.meas tran t_dis TRIG v(vp) val='vinit' FALL=1 TARG v(vp) val='vdd*0.25' FALL=1

.tran 1n 1.5m sweep DATA=input

.DATA input
+ vdd vinit
+ 0.400 0.120
+ 0.400 0.160
+ 0.400 0.200
+ 0.400 0.240
+ 0.400 0.280
+ 0.400 0.320
+ 0.400 0.360
+ 0.400 0.400
+ 0.450 0.135
+ 0.450 0.180
+ 0.450 0.225
+ 0.450 0.270
+ 0.450 0.315
+ 0.450 0.360
+ 0.450 0.405
+ 0.450 0.450
+ 0.500 0.150
+ 0.500 0.200
+ 0.500 0.250
+ 0.500 0.300
+ 0.500 0.350
+ 0.500 0.400
+ 0.500 0.450
+ 0.500 0.500
+ 0.550 0.165
+ 0.550 0.220
+ 0.550 0.275
+ 0.550 0.330
+ 0.550 0.385
+ 0.550 0.440
+ 0.550 0.495
+ 0.550 0.550
+ 0.600 0.180
+ 0.600 0.240
+ 0.600 0.300
+ 0.600 0.360
+ 0.600 0.420
+ 0.600 0.480
+ 0.600 0.540
+ 0.600 0.600
+ 0.650 0.195
+ 0.650 0.260
+ 0.650 0.325
+ 0.650 0.390
+ 0.650 0.455
+ 0.650 0.520
+ 0.650 0.585
+ 0.650 0.650
+ 0.700 0.210
+ 0.700 0.280
+ 0.700 0.350
+ 0.700 0.420
+ 0.700 0.490
+ 0.700 0.560
+ 0.700 0.630
+ 0.700 0.700
+ 0.750 0.225
+ 0.750 0.300
+ 0.750 0.375
+ 0.750 0.450
+ 0.750 0.525
+ 0.750 0.600
+ 0.750 0.675
+ 0.750 0.750
+ 0.800 0.240
+ 0.800 0.320
+ 0.800 0.400
+ 0.800 0.480
+ 0.800 0.560
+ 0.800 0.640
+ 0.800 0.720
+ 0.800 0.800
.ENDDATA
