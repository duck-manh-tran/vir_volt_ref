module da_mult (clk, rst_n, mult_dn, inst_a, inst_b, mult_out);

endmodule
